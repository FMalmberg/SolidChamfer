MZ�       ��  �       @                                   �   � �	�!�L�!This program cannot be run in DOS mode.
$       3�Q�w�?�w�?�w�?����v�?�ܡ�j�?�ܕ��?�~Ҭ�t�?�w�>�=�?�ܔ�8�?�ܤ�v�?�ܢ�v�?�Richw�?�                        PE  L �HR        � !
  �  �      D�     �                       �         @                   @ L   l (                            ` �&  P�                            h� @            �                           .text   �     �                   `.rdata  �a   �  b   �             @  @.data    4         �             @  �.reloc   5   `  6                @  B                                                                                                                                                                                                                                                                                                                                                                                        �p���� �����U��V���p��� �Et	V�C�  ����^]� ���������U��EVP���� �p���^]� ����U��M��3���tD�����?w��    P���  ����u(�MQ�M��E    �� hH��U�R�E�p���� ��]� �������U���L�M�U�E�P�EQ�MRP�B �MĉE����  �M����  �}� �E�    ��  SVW�U��E�3�V�M�Q���UQ�MR�N �Mȋ�M�3�3�I�uԉE؉]܉u��U�u����  ��$    �M�9M�u�U��}�B��U��M�U��Mč<�;�sd;�w`+���;�uL��+��������?�  ��+�A��;�v-�������?+�;�s3���;�s��R�M��+N  �]܋E؋uԅ�t_����X;�uL��+��������?��  ��+�A��;�v-�������?+�;�s3���;�s��R�M���M  �]܋E؋uԅ�t���Uċ}������E�;Mu�L�;Mt��;M��   �M9L���   �U��M����U;�sh��;�wb��+���;�uL��+��������?�  ��+�A��;�v-�������?+�;�s3���;�s��R�M��%M  �]܋E؋uԅ�t`����Y;�uL��+��������?��  ��+�A��;�v-�������?+�;�s3���;�s��R�M���L  �]܋E؋uԅ�t�M����E؋M��U�AJ�M�;�������M̋Uč|��;�sd;�w`+���;�uL��+��������?�(  ��+�A��;�v-�������?+�;�s3���;�s��R�M��AL  �]܋E؋uԅ�t_����X;�uL��+��������?��  ��+�A��;�v-�������?+�;�s3���;�s��R�M���K  �]܋E؋uԅ�t���UċM̋L�����E�;Mu�:;}t;M��   �M9
��   �UȋM����U;�se��;�w_��+���;�uI��+��������?�(  +ދ�A��;�v*�������?+�;�s3���;�s��P�M��AK  �E؋uԅ�t]����V;�uI��+��������?��   +ދ�A��;�v*�������?+�;�s3���;�s��P�M���J  �E؋uԅ�t�M����UȋM�RV+�Q��P�M�� �U��E���}�]j QW��� j �U�RW���� 3�;�t	V��  ���E�@�}ԉ}؉}܉E�;E������_^[�E��MPQ�M� �M��e �M��] ��]�hx��Ҷ ���������������U�����  ��u3���]���  ��t�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�эU�R�( ��5�H�A�U�R�Ѓ��   ��]�����������������U��EHt3�]ù�5�)L �����]�̋��@    �     Ë�������������̋A�������������U��U�V�u�;�u�B;F��^]� U��UV�u���M;�|�M�	�;�^�M|�M��P]� �̋�3ɉ�H�H�Hf�H�������������U��E;u�A]� �A]� ��������U��E;u
�U�Q]� �E�A]� ��U��E;u�A]� �A]� ��������U��E;u
�U�Q]� �E�A]� ��U��V�uW�}���M;�|�M�;�_�^�M|�M�	�H�P�Hf�@  ]� ����U��E�H�y) u����H�y) t�]����U��E��y) u������y) t�]�����U��U�BV�0�r�0�~) u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~) u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ��������̋���z) u@�J�y) u��z) u��I �ʋ�z) t��ËR�z) u�;Ju��R�z) t������̋���y) t�I�Ë�z) u�J�y) u0�ыJ�y) t��ËQ�z) u�;
u��R�z) t��y) u��������������U��SVW���G�p�~) ��u$�EP�NQ���������t�v��ދ6�~) tދ�_^[]� ���������������U��A=H�$	r�EP��  ��h��蠲 @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z(��  V��    �P�r;��   �v8^(u�B(�F(�P�R�Z(�@�@�Q  ;Bu:�P�2�p�28^)u�F�p�r�q;Fu�V��p;u���V��P�P�B(�P�R�Z(�P�R�2�~�:�~8_)u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^(u�B(�F(�P�R�Z(�@�@�   ;u<��r�0�r8^)u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B(�P�R�Z(�P�R�r�>�z�>8_)u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z(�q���^�A�H�E�8_�A([]� �����������U��M��t+�E���P�Q�P�Q�P�Q�P�Q�P�Q�@�A]����������U��QSVW���G�p�~) �M�ذ�E�u@��} �A�ދ�tP�FP�)��������
�VRP�����E���t�6��v�~) �Mt���u��t8�G;u#QSj�MQ��������E_^��@[��]� �M�F����u�M�AP�FP��������t(�M�U�QSR�EP���������E_^��@[��]� �UR�\�  �E��_�0^�@ [��]� �������U��j�h��d�    P��SVW�`#3�P�E�d�    �e���j,��  �����u�3�;�t^�O��W�V�O�Nf�F(�E��UR�FP��W�U������E������ƋM�d�    Y_^[��]� �M�Q��  ��3�PP�ݰ �E�UR�M��ʯ �E�p�hH��E�P蹰 ������������U����ESVW��M�^PQ�M�������W���H����E;Ft%��PW���T�����u�E� _3�;�^��[��]� �V�E�U� _3�;�^��[��]� U���0S�]VW�}W��S�M��������P�M�H�U�P�@W�M�S�M��U��E������P���f  �M�U��M�P�U��H�M�_^�P�H[��]� U���S�]VW��M�FSQ�M��E�������W���e����E;Ft��PW���q�����u�E�	�V�U��E��M�9u�USR���,����ESP�M��_���P����  _^[��]� ��������������U���SV��~ �FW�}�_uW�}PjW�)�����_^[��]� �M;u1��QS����������>  �MW�}QjW���������_^[��]� ;�u7�@��SP���������  �V�BW�}Pj W��������_^[��]� ��QS���o�����t^�M�M�M������US��R���N�����t=�E�H�y) W�}��tPj W�_�����_^[��]� �URjW�H�����_^[��]� �ES��P���������te�M�M�M�����E;Ft��PS���������t?�E�M�Q�z) W�}tQj W���������_^[��]� PjW���������_^[��]� j W�E�P���'�����E_^�[��]� �������U���0SVW�}W���<�����;^t�CPW���I�����tW�M�������W�MЋ�M؋H�UԋP�M��U܋P�@�M�Q�ΉU�E�����PS�UR��������E_^��[��]� _^�C[��]� �̡�5�PH���   h�  Q�Ѓ�������̡�5�PH���   h�  Q�Ѓ��������U��VW�����5�QHh�  P���   �Ћu��;�}*��5�?�QH���   j h�  W�Ѓ��v_��^]� ��5��JH���   h�  P�ҋO��+��v_��^]� ���������������U��V����5�QHWh�  P���   �Ћ}��5�QH��;�} �6���   j h�  V�Ѓ����_^]� �h�  P���   �Ћȋǃ�+���F_^]� ��������U���3ɉH�H�H�H�H�H�M�]� ��������������U���SV����5�QHWh�  P���   �Ћ�5�QH�؋h�  P���   �ЋN+N�����Q�N+N�E�����*����������P�.I ���5�QHj h�  P���   �Ћ�5�QH�E��j h�  P���   �ЋN+N�E�����*����������3��td�M��[3ҍ��
��$    �U��F��X�Y�X�Y�X�Y�X�Y�@�A���U��V+V����*��������G�;�r��N+N3�����tA�M���3�M�    �F��X�Y�X�Y�@�A�F+FG������;�rЋN�V;�t5��;�t,�8�9�x�y�x�y�x�y�x�y�x�y����;�uԉN�N�V;�t*��;�t!��8�9�x�y�x�y�x�y����;�u��N_^[��]�������U��VW���EP�O�M  �O+O�?����*���5�������QH���   h�  W�Ѓ�_�D0�^]� U��S�ًC�MVW;�s?�K�U;�w5��+�;Cu
j�K�  �C���{��tB���W�P�O�H�W�*;Cu
j�K�P  �C��t�M��U�P�M�H�U�P�C�{���5+{�QHh�  P���   ���Ѓ��D8�_^[]� ��������������U��M��3���tF�����
w�I���P�
�  ����u(�MQ�M��E    �)� hH��U�R�E�p��� ��]� �����U��M��3���t@�����w��Q��  ����u(�EP�M��E    �Ϧ hH��M�Q�E�p�辧 ��]� �����������U��E��t%�M���Q�P�Q�P�Q�P�Q�P�I�H]����������������U��E��t�M���Q�P�Q�P�I�H]������������U��j�hТd�    PQSVW�`#3�P�E�d�    �e��E�    �]�}�u��$    ;utVWS�C��������}���u���E������ǋM�d�    Y_^[��]�j j 軦 ��������������U��j�h�d�    PQSVW�`#3�P�E�d�    �e��E�    �]�}�u��$    ;utVWS����������}���u���E������ǋM�d�    Y_^[��]�j j �+� ��������������U��E�UP�Ej ��Q�MQRP�������]� �����������U��E�UP�Ej ��Q�MQRP�"�����]� �����������U��j�h�d�    P��SVW�`#3�P�E�d�    �e���}�����
v
hx��Q� �N+����*���������;�shW�N������E��E�    P�NQ�R���"����E�������N+˸���*�����������t	S���  ���E�@�E�ȉV��ȉV��M�d�    Y_^[��]� �E�P��  ��j j �Ф ���U��j�h0�d�    PQSVW�`#3�P�E�d�    �e���]�����v
hx��c� �F+��;�sRS�N�k����E�E�    P�NQ�R���r����E�������~+���t	P�
�  �����E؉^�����~��M�d�    Y_^[��]� �EP���  ��j j �� ���������U��QVW�9+׸���*��E������򺪪�
+�;�s
hx�螡 �Q�+׸���*���������;�v!���꿪��
+�;�s3���;�s��P�����_^]� ��������U��A�UV�1W+ƿ�����+�;�s
hx��,� Q+���;�v!�������+�;�s3���;�s��R�Z���_^]� ����U��V�uW���O;�sb�;�w\+𸫪�*���������;Ou	j���������v���G��tc���Q�P�Q�P�Q�P�Q�P�I�H�G_^]� ;Ou	j�������G��t"���N�H�V�P�N�H�V�P�N�H�G_^]� ������������U��E�H�y u����H�y t�]���̋A�������������U��QV��EP�M�Q���j  �3�;V^����]� ���������U���Vj �EP���l  P�M�Q���;  ^��]� ���������U��U�BV�0�r�0�~ u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~ u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ��������̋���y t�I�Ë�z u�J�y u0�ыJ�y t��ËQ�z u�;
u��R�z t��y u��������������U��A=���?r�EP�Z�  ��h���`� @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z��  V��    �P�r;��   �v8^u�B�F�P�R�Z�@�@�Q  ;Bu:�P�2�p�28^u�F�p�r�q;Fu�V��p;u���V��P�P�B�P�R�Z�P�R�2�~�:�~8_u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^u�B�F�P�R�Z�@�@�   ;u<��r�0�r8^u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B�P�R�Z�P�R�r�>�z�>8_u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z�q���^�A�H�E�8_�A[]� �����������U��j�hP�d�    P��SVW�`#3�P�E�d�    �e���j��  �����u�3�;�t^�O��W�V�O�Nf�F�E��UR�FP��W蕱  ���E������ƋM�d�    Y_^[��]� �M�Q��  ��3�PP�ݝ �E�UR�M��ʜ �E�p�hH��E�P蹝 ������������U��Q�Q�B�x W�}uV�79p}�@��Ћ �x t�^�A�U;�t�;J|�E��E�_��]� �E��E���E�_��]� ��������������U�����E��������u����]��ر������u
���б]�]�x� ��������U��V�u�F��F�����������������\� ��������������D�Ez��^�P�P�]��������������N�X�N^�X]���������������U�조5�E�P�E���   ���$P��]� �����������̡�5�P@�B,Q�Ѓ����������������U�조5�PH�EP�EPQ���   �у�]� ������������̡�5�PH��p  j h�  Q�Ѓ�����̡�5�PH��p  j h�  Q�Ѓ������U��M�Q���VW�y�I;׍I�Ru3�u�֍֍@�$ƍ��B���`�B�`�� �A�`�A�`�8�4@�E�Ѝ��$��4��B�f�B��f���ȍ��"�@�b�@�b���u�̍U���R��V���]������������]��������]�������_��^��]�����������U�조5�Pl�E�I�RPQ�҃�]� �U��V�u��tIS�]W�}VW���$A ��5���   �B4����PWS�������5���   �B(�����Ћ���u�_[^]����������U�조5�H@�U�A,VR������5�QQ���$�B,h�  ���Ћ�5�Q�B4j h�  ���Ћ�5�Q�B4h�  h�  ���и   ^]� ���������������U�조5�H�A��4�U�VR�Ћ�5�Q�Jj j��E�h�P�ы�5�B�P�M�Q�ҡ�5�H�Aj j��U�h��R�Ћ�5�Q�J�E�P�ы�5�B�Pj j��M�hܲQ�҃�<�E�P�M��] � j P�M�Qh`> j�U�Rh[� �h ���M����^ ��5�H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�P�M�Q�҃���^��]������������U����   SVW�}����> ��5���   �B4���Ћ�3�;�uVV�G ��_^[��]� ��5�u��u��u��uĉuȉuЉű��   �BT���ЍM�Qh�   �E��]���	 ����u�M��� _^3�[��]� ��5���   �MЋ��   V�ҋ�5���   �Bh�  ���Ѕ�uPP��F ���M����~ _��^[��]� �MSQ���W> ��5���   �P4����P�EPW�����������= ���> ��5�Q@�B,W�Ћ؃��]���^ ��5�E�Q���   j h�  ���Ћ�5�QH�؋��   h�  V�Ћ�5�QHj �E􋂘   h�  V�Ѝ���������Z  �$�L; �MQ���4 �<  �M��~J�   �X�M�M�W�R�^ �M�G�P�^ �MW�^ �;Kt�M�WR�^ �����Mu��EP���5 ��  j h�  ����������  ���S�����5�Q�����   j h�  ���Ѕ���  ��5�Q���   3�Sh�  ���Ѕ�t�MQ���%4 ����^ ����$��h�  �����]��M��= S���W���P���?���P���'���P�M��.= �]9]���   �]�������E���P�����P��,���R� ���� �]����@�M��]��@�EP�]��������3��<��th������������P������P�����R������ �@���@���M����M������M����$�<����E���������Az�E��Q�M��\ G��|��E�E�@�E;E��5����UR����3 �M��!< �A��5���   �BT���Ћ�5�Q�M�j P�Blh�  �Ѕ�t�MQ����e ���~] 3�jP�]�袼  ��;��O  �E؉ �E؉@�E؉@�U��BH�E�V��D����@I�,  �ES��D���Q�U�RPV��  ��5�Q�M����   ��Sh�  �����5�Q�M����$�����   h�  ���]�;�~�M�Q��D����=  Ou��(�  SV�ȉE���  �E�U����$RV�M���  ��5�HH���   jV�ҋM���SSS���  ��5���   �BSj���ЍM�Q���  ����D����]��  �E؋PQ�UR�M��  �E�P�j�  �MQ��Z ���M��]� _��^[��]� �UR�M�]�r� hH��E�P�E�p��a� o7 �9 7 �7 ����U��U�V�p�2�p�~I u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��E�H�yI u����H�yI t�]����U��E��yI u������yI t�]�����U��U�V�p�2�p�~ u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��E��y u������y t�]����̋���zI u@�J�yI u��zI u��I �ʋ�zI t��ËR�zI u�;Ju��R�zI t������̋���z u@�J�y u��z u��I �ʋ�z t��ËR�z u�;Ju��R�z t������̋���z u@�J�y u��z u��I �ʋ�z t��ËR�z u�;Ju��R�z t�������U��U�BV�0�r�0�~I u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��U�BV�0�r�0�~ u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��V���UR �Et	V�)�  ����^]� ���������������Vh��jh�5j輺  ������t����Q �����^�3�^���������������U���S�]�{I VW�M�t
h ��� �M�]�������yI t�{��C�xI t���
�E�x;�ur�I �su�w�M��A9Xu�x�9u�>��~�A9u�I t���W�����M����Q��I�M�9Yux�I t�ƉA�kW�k����M���A�Z�A��;Cu����I �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�SH�HH�PH�KH�E��8XH��   �M��Q;z��   8_H��   �;�ue�F�xH u�XHV�FH �t����F�M��xI ut�8ZHu�P8ZHta�P8ZHu��ZHP�@H �2����F�M��VH�PH�^H�@V�XH�'����t�xH u�XHV�FH ������M��xI u�P8ZHu�8ZHu�@H �A���v;x�J����0�8ZHu�P�ZHP�@H �������M��VH�PH�^H� V�XH�����_H�M�Q襷  �M��A��_^[��tH�A�E�U���]� ���U���S�]�{ VW�M�t
h ���� �M�]�������y t�{��C�x t���
�E�x;�ur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W�4�  �M����Q��I�M�9Yux� t�ƉA�kW�����M���A�Z�A��;Cu���� �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S�H�P�K�E��8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F �����F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ ������F�M��V�P�^�@V�X�G����t�x u�XV�F ������M��x u�P8Zu�8Zu�@ �A���v;x�J����0�8Zu�P�ZP�@ �������M��V�P�^� V�X�1����_�M�Q�U�  �M��A��_^[��tH�A�E�U���]� ���U���S�]�{ VW�M�t
h ��q� �M�]�������y t�{��C�x t���
�E�x;�ur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W�����M����Q��I�M�9Yux� t�ƉA�kW�  �M���A�Z�A��;Cu���� �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S�H�P�K�E��8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F �4����F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �2����F�M��V�P�^�@V�X������t�x u�XV�F ������M��x u�P8Zu�8Zu�@ �A���v;x�J����0�8Zu�P�ZP�@ ������M��V�P�^� V�X�����_�M�Q��  �M��A��_^[��tH�A�E�U���]� ���U��SVW�}�I �ً�u�FP��������6W躲  ���~I ��t�_^[]� ��������U��SVW�}� �ً�u�FP��������6W�z�  ���~ ��t�_^[]� ��������SVW���G�X�{I ��u�NQ���b����6S�:�  ���~I ��t�G�@�G� �G�@�G    _^[����SVW���G�X�{ ��u�NQ���r!  �6S��  ���~ ��t�G�@�G� �G�@�G    _^[����U��Q�UV��F�M;u;�u���A����F��E�^��]� ;�t^�yI ��uB�A�xI u�ȋ�xI u��ȋ�xI t��M��A�xI u;Hu�ȉM�@�xI t�ER�U�R���f����M;Mu��E�^��]� ��U��Q�UV��F�M;u;�u����  �F��E�^��]� ;�t^�y ��uB�A�x u�ȋ�x u��ȋ�x t��M��A�x u;Hu�ȉM�@�x t�ER�U�R�������M;Mu��E�^��]� ��U��Q�UV��F�M;u;�u���Q����F��E�^��]� ;�t^�y ��uB�A�x u�ȋ�x u��ȋ�x t��M��A�x u;Hu�ȉM�@�x t�ER�U�R��������M;Mu��E�^��]� ��U��QV��FH�WPQ�E�P�N@�E����NHQ輯  �F4���PQ�U�R�N0�����F4P蝯  �F$���PQ�M�Q�N �g����V$R�~�  �F3���;�t	P�l�  ���~�~�~�;�t	P�T�  ���>�~�~_^��]����U���SV��W3��>�~�~�~�~�~j�~(��  ��;���   �F$� �F$�@�F$�@�F$��X�N$�Yj�~8��  ��;���   �F4� �F4�@�F4�@�V4�Z�F4�M��X������@j�N@�FD�~L蟬  ��;�t.�FH� �FH�@�FH�@�NH�E�Y�VH�Z�FT_��^[��]� �MQ�M�}蔃 hH��U�R�E�p�胄 �EP�M�}�p� hH��M�Q�E�p��_� �UR�M�}�L� hH��E�P�E�p��;� ��������������U���V��jP�F    �٫  ����t&�F� �F�@�F�@�N��AH�V�BI��^��]ÍE�P�M��E�    �҂ hH��M�Q�E�p���� ���̋���yI t�I�Ë�zI u�J�yI u0�ыJ�yI t��ËQ�zI u�;
u��R�zI t��yI u��������������U��A=#I�r�EP�
�  ��h���� @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8ZH��  V��    �P�r;��   �v8^Hu�BH�FH�P�R�ZH�@�@�Q  ;Bu:�P�2�p�28^Iu�F�p�r�q;Fu�V��p;u���V��P�P�BH�P�R�ZH�P�R�2�~�:�~8_Iu�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^Hu�BH�FH�P�R�ZH�@�@�   ;u<��r�0�r8^Iu�F�p�r�q;Fu�V��p;Fu�V���B�P�P�BH�P�R�ZH�P�R�r�>�z�>8_Iu�W�z�~�y;Wu�w��z;u�7��w��}�r�P8ZH�q���^�A�H�E�8_�AH[]� �����������U��Q�US�ًK�A�xI V��W�M�u-�z�} ��t9x���;x���M���t� ��@�xI t֋��}��t5�C�M;0u RVjQ���e�����E_^��@[��]� ������}�U�GR;B}$�M�VQ�UR���-�����E_^��@[��]� �4�  �E���8_^�@ [��]� ���������������U��E��t�M�VW�q�x�   ��_^]�������������U�조5��SVW�}j �ًHH���   h�  W�ҋC�0��;���   �E�N�F0j �ɍE��F8P��Q�F@�M��W�F�����]��F �]��F(�]��O�  �~I u@�F�xI u����xI u-��    ����xI t���F�xI u;pu���@�xI t���;s�v������0 _^[��]� U��VW�EP�  �   �u���_^]�4 U��VW�EP�  ���E�   ���_^]� ��������������U���V��~ �FW�}uW�}PjW�}�����_^��]� S�];u&�O;K��   W�}SjW���P���[��_^��]� ;�u'�@�P;W��   W�}Pj W�%���[��_^��]� �G;C}M�M�]�����E�O9H}7�H�yI W�}��tPj W�����[��_^��]� SjW�����[��_^��]� �G9C}R�M�]������E;Ft�O;H}7�S�zI W�}��tSj W����[��_^��]� PjW�v���[��_^��]� j W�E�P��������E[_�^��]� �������������U��U��8VW���O�A�xI ��u�
�I 9H}�@���� �xI t�;wt�;F}M��
���U����M���R�Ë������]����]��]��]��]��]��nE  PV�EP���!����E_��^��]� _�F^��]� ��������U����U���P�M�P��P(�P �X��M�P�U�H�M�P�U�H�M �H�M(�P�U$�P�U,�H �M0�P$�U4�H(�P,]�0 �������������U��E�H�y u����H�y t�]����U��E��y u������y t�]�����U��E��y! u������y! t�]�����U��E�H�y u����H�y t�]���̋���z u@�J�y u��z u��I �ʋ�z t��ËR�z u�;Ju��R�z t������̋���y t�I�Ë�z u�J�y u0�ыJ�y t��ËQ�z u�;
u��R�z t��y u�������������̋���y t�I�Ë�z u�J�y u0�ыJ�y t��ËQ�z u�;
u��R�z t��y u�������������̋���z! u@�J�y! u��z! u��I �ʋ�z! t��ËR�z! u�;Ju��R�z! t�������U��U�BV�0�r�0�~ u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~ u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��U�BV�0�r�0�~ u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��U�V�p�2�p�~ u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��U�BV�0�r�0�~! u�V�r�p�I^;Qu�A��B]� �J;u���B]� �A��B]� �������������U��SVW���G�p�~ ��u$�EP�NQ��������t�v��ދ6�~ tދ�_^[]� ���������������U��M�E+�V���4�    �EVQP�x ���^]� �����U��A=���r�EP���  ��h��� v @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z��  V��    �P�r;��   �v8^u�B�F�P�R�Z�@�@�Q  ;Bu:�P�2�p�28^u�F�p�r�q;Fu�V��p;u���V��P�P�B�P�R�Z�P�R�2�~�:�~8_u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^u�B�F�P�R�Z�@�@�   ;u<��r�0�r8^u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B�P�R�Z�P�R�r�>�z�>8_u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z�q���^�A�H�E�8_�A[]� �����������U��A=���r�EP�ʟ  ��h����s @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z ��  V��    �P�r;��   �v8^ u�B �F �P�R�Z �@�@�Q  ;Bu:�P�2�p�28^!u�F�p�r�q;Fu�V��p;u���V��P�P�B �P�R�Z �P�R�2�~�:�~8_!u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^ u�B �F �P�R�Z �@�@�   ;u<��r�0�r8^!u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B �P�R�Z �P�R�r�>�z�>8_!u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z �q���^�A�H�E�8_�A []� �����������U��A=TUUr�EP蚝  ��h���q @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z��  V��    �P�r;��   �v8^u�B�F�P�R�Z�@�@�Q  ;Bu:�P�2�p�28^u�F�p�r�q;Fu�V��p;u���V��P�P�B�P�R�Z�P�R�2�~�:�~8_u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^u�B�F�P�R�Z�@�@�   ;u<��r�0�r8^u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B�P�R�Z�P�R�r�>�z�>8_u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z�q���^�A�H�E�8_�A[]� �����������U��A=���r�EP�j�  ��h���po @S�A�EW�}�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z��  V��    �P�r;��   �v8^u�B�F�P�R�Z�@�@�Q  ;Bu:�P�2�p�28^u�F�p�r�q;Fu�V��p;u���V��P�P�B�P�R�Z�P�R�2�~�:�~8_u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^u�B�F�P�R�Z�@�@�   ;u<��r�0�r8^u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B�P�R�Z�P�R�r�>�z�>8_u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z�q���^�A�H�E�8_�A[]� �����������U��j�hp�d�    P��SVW�`#3�P�E�d�    �e���j��  �����u�3�;�t^�O��W�V�O�Nf�F�E��UR�FP��W��  ���E������ƋM�d�    Y_^[��]� �M�Q輘  ��3�PP��n �E�UR�M���m �E�p�hH��E�P��n ������������U��j�h��d�    P��SVW�`#3�P�E�d�    �e���E=���?v
hx��Rl �N+��;�sSP�N�����؉]��E�    S�VR�P��������E�������~+�����t	P���  ���M���V���F��M�d�    Y_^[��]� �M�Q�×  ��j j ��m �������U���S�]�{ VW�M�t
h ���k �M�]�������y t�{��C�x t���
�E�x;�ur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W������M����Q��I�M�9Yux� t�ƉA�kW�����M���A�Z�A��;Cu���� �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S�H�P�K�E��8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F ������F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �����F�M��V�P�^�@V�X�����t�x u�XV�F �������M��x u�P8Zu�8Zu�@ �A���v;x�J����0�8Zu�P�ZP�@ �:�����M��V�P�^� V�X�����_�M�Q腕  �M��A��_^[��tH�A�E�U���]� ���U���S�]�{ VW�M�t
h ��i �M�]��������y t�{��C�x t���
�E�x;�ur� �su�w�M��A9Xu�x�9u�>��~�A9u� t���W������M����Q��I�M�9Yux� t�ƉA�kW�����M���A�Z�A��;Cu���� �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S�H�P�K�E��8X��   �M��Q;z��   8_��   �;�ue�F�x u�XV�F �T����F�M��x ut�8Zu�P8Zta�P8Zu��ZP�@ �����F�M��V�P�^�@V�X�����t�x u�XV�F �R�����M��x u�P8Zu�8Zu�@ �A���v;x�J����0�8Zu�P�ZP�@ ������M��V�P�^� V�X������_�M�Q�5�  �M��A��_^[��tH�A�E�U���]� ���U���S�]�{! VW�M�t
h ��Qg �M�]��&�����y! t�{��C�x! t���
�E�x;�ur�! �su�w�M��A9Xu�x�9u�>��~�A9u�! t���W�t����M����Q��I�M�9Yux�! t�ƉA�kW�z  �M���A�Z�A��;Cu����! �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S �H �P �K �E��8X ��   �M��Q;z��   8_ ��   �;�ue�F�x  u�X V�F  ������F�M��x! ut�8Z u�P8Z ta�P8Z u��Z P�@  ��z  �F�M��V �P �^ �@V�X �w����t�x  u�X V�F  �z  ��M��x! u�P8Z u�8Z u�@  �A���v;x�J����0�8Z u�P�Z P�@  ������M��V �P �^ � V�X �1z  �_ �M�Q��  �M��A��_^[��tH�A�E�U���]� ���U��SVW�}� �ً�u�FP��������6W蚐  ���~ ��t�_^[]� ��������U��SVW�}� �ً�u�FP��������6W�Z�  ���~ ��t�_^[]� ��������U��SVW�}�! �ً�u�FP��������6W��  ���~! ��t�_^[]� ��������U��Q�US�ًK�A�x V��W�M�u-�z�} ��t9x���;x���M���t� ��@�x t֋��}��t5�C�M;0u RVjQ���%�����E_^��@[��]� �����}�U�GR;B}$�M�VQ�UR���������E_^��@[��]� �D�  �E���8_^�@ [��]� ���������������U��QSVW���G�p�~ �M�ذ�E�u@��} �A�ދ�tP�FP�	��������
�VRP������E���t�6��v�~ �Mt���u��t8�G;u#QSj�MQ��������E_^��@[��]� �M�f����u�M�AP�FP��葬����t(�M�U�QSR�EP���I�����E_^��@[��]� �UR�<�  �E��_�0^�@ [��]� �������U��Q�US�ًK�A�x! V��W�M�u-�z�} ��t9x���;x���M���t� ��@�x! t֋��}��t5�C�M;0u RVjQ���������E_^��@[��]� �v  �}�U�GR;B}$�M�VQ�UR��������E_^��@[��]� �d�  �E���8_^�@ [��]� ���������������U��QSVW���G�p�~ �M�ذ�E�u@��} �A�ދ�tP�FP�)��������
�VRP�����E���t�6��v�~ �Mt���u��t8�G;u#QSj�MQ��������E_^��@[��]� �M�&����u�M�AP�FP��豪����t(�M�U�QSR�EP���������E_^��@[��]� �UR�\�  �E��_�0^�@ [��]� �������U��Q�US�ًK�A�x V��W�M�u-�z�} ��t9x���;x���M���t� ��@�x t֋��}��t5�C�M;0u RVjQ���U�����E_^��@[��]� �����}�U�GR;B}$�M�VQ�UR��������E_^��@[��]� 脋  �E���8_^�@ [��]� ���������������U��A�UV�1W+ƿ���?��+�;�s
hx��L_ Q+���;�v!�������?+�;�s3���;�s��R����_^]� ����U��j�h��d�    P��SVW�`#3�P�E�d�    �e��ى]�C�E�}� uO�OQ���f������U�V�G�F�M�y t�u��E�    V�R�������V�GP���|����F�E������E�M�d�    Y_^[��]� �M�Q�M������j j �` ������SVW���G�X�{ ��u�NQ���b����6S��  ���~ ��t�G�@�G� �G�@�G    _^[����SVW���G�X�{ ��u�NQ���R����6S�ʉ  ���~ ��t�G�@�G� �G�@�G    _^[����SVW���G�X�{! ��u�NQ���B����6S�z�  ���~! ��t�G�@�G� �G�@�G    _^[����U���V��~ �FW�}uW�}PjW�M�����_^��]� S�];u&�O;K��   W�}SjW��� ���[��_^��]� ;�u'�@�P;W��   W�}Pj W�����[��_^��]� �G;C}M�M�]�7q  �E�O9H}7�H�y! W�}��tPj W����[��_^��]� SjW����[��_^��]� �G9C}R�M�]�����E;Ft�O;H}7�S�z! W�}��tSj W�Z���[��_^��]� PjW�F���[��_^��]� j W�E�P���������E[_�^��]� �������������U���SV��~ �FW�}�_uW�}PjW������_^[��]� �M;u1��QS���˥�����>  �MW�}QjW���������_^[��]� ;�u7�@��SP��蓥�����  �V�BW�}Pj W��������_^[��]� ��QS���_�����t^�M�M�M�����US��R���>�����t=�E�H�y W�}��tPj W�O�����_^[��]� �URjW�8�����_^[��]� �ES��P��������te�M�M�M������E;Ft��PS���Ȥ����t?�E�M�Q�z W�}tQj W���������_^[��]� PjW���������_^[��]� j W�E�P��������E_^�[��]� �������U���V��~ �FW�}uW�}PjW������_^��]� S�];u&�O;K��   W�}SjW���p���[��_^��]� ;�u'�@�P;W��   W�}Pj W�E���[��_^��]� �G;C}M�M�]�����E�O9H}7�H�y W�}��tPj W����[��_^��]� SjW�����[��_^��]� �G9C}R�M�]�����E;Ft�O;H}7�S�z W�}��tSj W����[��_^��]� PjW����[��_^��]� j W�E�P��������E[_�^��]� �������������U��j�hУd�    P��SVW�`#3�P�E�d�    �e���j謂  �����u�3�;�t^�O��W�V�O�Nf�F�E��UR�FP��W�n  ���E������ƋM�d�    Y_^[��]� �M�Q�L�  ��3�PP�}Z �E�UR�M��jY �E�p�hH��E�P�YZ ������������U��E��t�M���A�X]��������U��E��t�M���I�H]��������U�����PS�ك{ ��   �C�U�V�U�0�U��U�;���   W�}������؋F��P�M�Q�������@�~! �E��U��@ �E��U��@(�E��U��F�E��U�u:�F�x! u����x! u'����x! t���F�x! u;pu���@�x! t���;su���_������������D{%�؋E��^��[������������X���X��]� �������؋E�P^�P[���]� �E�[�P�X��]� �������U���V�q@j �EP���I���P�M�Q���m���^��]� ������U���V�q j �EP���)���P�M�Q���]���^��]� ������U���V�q0j �EP�������P�M�Q���-���^��]� ������U��QV��EP�M�Q�N 虺���3�;V$^����]� ��������U��QV��EP�M�Q�N0�i����3�;V4^����]� ��������U��EP�d  ]� U��EP���Q  ]� �������������U���   �ESV�uWVP�M�负���}��S��������E�;Gt��PS���s�����u�E��	�O�M��E�� ;Gt�@_^[��]� ��M������������X�X�ѭ���U�]��R�E�P������� �]�V�@�M��]�Q�@���]�������U��R��x���P��������F�@��0�@ ���F �@(���F(W�@��������E��E��E�����X�X���X�X �X(�s����M�UQR�M�賞���MP�Z!  �8��_^[��]� �������������U���  SVW3�j$��}��6~  ��;���  �E�� �E��@�E��@�E��@ �M��A!�VTR��@���荪���~�^+>+^�FT��5�QHj h�  P���   �����}��]��Ѓ��M��E�謝����M��Pj�U��E�    �}  3Ƀ�;���  �E�� �E��@�E��@�E��@�U��Bj��$����j}  3Ƀ�;���  �� ���� �� ����@�� ����@�� ����@�� ����B�M�;���  �d$ ��M̋��E����<�\�LP�M�M��@���PQ�U܍U�RSW�Ή}�]��N����M�E���@���P�E�Q�M�U�RPQ���-����V$�ʉE�A�x u9x}�@��ȋ �x t�F$�M�;�t
;y|�E���EЍE�9u?�U��E�P�M��U��.  �M�Q���=!  ��U��R�M��}���-  �M�Q���!  ����V$�ʋA�x u9X}�@��ȋ �x t�F$�M�;�t
;Y|�E���E؍E�9u?�U��E�P�M��U��-  �M�Q���   ��U��R�M��]��k-  �M�Q���   ����~$�U�ϋA�x u9P}�@��ȋ �x t�F$�M�;�t
;Q|�E���E��E�98uB�U�E�P�M��U��-  �M�Q���<   ��U���E�P�M��U���,  �M�Q���   ����~$�U܋ϋA�x u��    9P}�@��ȋ �x t�F$�M�;�t
;Q|�E����d�����d���98uB�U�E�P�M��U��v,  �M�Q���  ��U���E�P�M��U��U,  �M�Q���  �����]̋���E�����P�ĉ�M��H�M�H��@����P肩���EԋF�U�;�sg��M�;�w^���N+���;�u@+���=���?�x  +�@��;�v&�������?+�;�s3���;�s��Q�������]̋F��t[�����R�N;�u?�+���=���?�  +�@��;�v#�������?+�;�s3���;�s��Q���8����F��t�Uԉ�F����U��E�ɉȋ���M�C҉L��]�;]��]����]�3ɉM�;���
  �V�Eԋ��]��E���P�M�H�@�U��M�E�;��>  ��@���P�E�S�M�QRP��������@���Q�M�S�U��E��E�RPQ���v����M荕@���R�U�S�E�E�PQR���X����V4�ʉE؋A�x u%�]�d$ 9X}�@�hx���N �ȋ �x t�F4�M�;�t�]�;Y|�E����d�����d����]�9tb�N4�A�x u9X}�@��ȋ �x t�F4�M�;�t
;Y|�E���E��E�9t$�E�j �M�Q�N0�E������P��L���R�N0�&����V4�ʋA�x u9X}�@��ȋ �x t�F4�M�;�t
;Y|�E���E�E�]�9to�N4�A�x u��$    9X}�@��ȋ �x t�F4�M�;�t
;Y|�E������������9t$�E�j �M�Q�N0�E��D���P��<���R�N0�t����V4�ʋA�x u��    9X}�@��ȋ �x t�F4�M�;�t
;Y|�E��������������9tk�N4�A�x �]�u9X}�@��ȋ �x t�F4�M�;�t
;Y|�E��������������9t$�E�j �M�Q�N0�E�荰��P��D���R�N0���������������@�������X�X�]����Mԋ؋F���E�P������]ЉU���  �M��]Q�����R���v���� ݝt���������@ݝ|����@�E�P�]�Q���M����U�M��R��|���P�8����@�C�M�Q������ݝ`���R�C �@ ݝh����C(�]�@(��ݝp��������݅`�����0�@�@ ܅h����@(��܅p����P�������݅t���݅|����E�����X���X���X�X �X(�E�P�����V4�]��ʋA�x u�I 9X}�@��ȋ �x t�F4�M�;�t
;Y|�E������������9u?�MЍU��M�R�M���&  �M�Q���  ��U��R�M��]��&  �M�Q����  ����V4�]�ʋA�x u9X}�@��ȋ �x t�F4�M�;�t
;Y|�E��������������9u?�UЍE�P�M��U��N&  �M�Q���  ��U��R�M��]��0&  �M�Q���e  ����^4�U؋ˋA�x u9P}�@��ȋ �x t�F4�M�;�t
;Q|�E���E��E�9�G  �UЍE�P�M��U���%  �M�Q����  ��U���E�P�M��U��%  �M�Q�   �M���@���R�U�S�E�PQR���S����U�E���@���P�E�S�M�QRP���5�����@���Q�M�S�U��E�E�RPQ�������M荕@���R�U�S�E؍E�PQR��������^4�ˉE̋A�x u�U���I 9P}�@��ȋ �x t�F4�M�;�t�U�;Q|�E���E��E�9tA�E��M�Q��T���R�N0�E�貭��9t$�E�j �M�Q�N0�E��ʬ��P��X���R�N0������E��M�Q��x���R�N0�E��q����^49tA�E�M�Q������R�N0�E��Q���9t$�E�j �M�Q�N0�E��i���P��|���R�N0�����E�M�Q������R�N0�E������^49tA�E܍M�Q������R�N0�E�����9t$�E�j �M�Q�N0�E�����P������R�N0�8����E܍M�Q������R�N0�E�诬���^49tA�E�M�Q������R�N0�E�菬��9t$�E�j �M�Q�N0�E�觫��P��l���R�N0����������������@�������X�X�w����Mԋ؋F���E�P������]ЉU���  �M��]Q������R������� ݝt����������@ݝ|����@�E�P�]�Q���g����U�M��R��|���P�R����@�C�M�Q�����ݝ����R�C �@ ݝ�����C(�]�@(��ݝ���������@������܅����ݝ�����@ ܅����ݝ�����@(�E�܅����PQ��ݝ����������@܅�����@ �U�܅������0�@(��܅����R�H���������݅t���݅|����E�����X�X���X�X �X(�_����E��M�Q������R�N0�E������ �]�;F4u?�M�Q�M��]���!  �U�R���  ��M���E�Q�M��E��!  �U�R����  ����E�M�Q�� ���R�N0�E�脪��� ;F4u?�M�Q�M��]��~!  �U�R���  ��M���E�Q�M��E��]!  �U�R���  ����E؍M�Q������R�N0�E��%���� ;F4u?�M�Q�M��]��!  �U�R���T  ��M���E�Q�M��E���   �U�R���3  ����E̍M�Q�U�R�N0�E��ɩ��� ;F4u?�M�Q�M��]���   �U�R����  ��M���E�Q�M��E��   �U�R����  ����E�@�E�;E��v����]S������  �E��8�}�;���   �d$ �GP������Q������� ݝt���������@Rݝ|����O�@������P�]�����݅t����݅|����P�E��������ʋH�������P�������H�������P��0����������������X���X݅�����X݅�����X ݅�����X(�GP������M��@����}ԋE�;��2����HQ�M���  �E��@�E�� �E�3ۉ@�]�9]���  ��$    �V����E��H�8�P�@;ȉE܍�@���P�M�MQ�U��E��U�RP�}��W��  ������U��@���Q�M�R�U��E��E�PQR��������M�E䍅@���P�E�Q�U�RWP�������N���E؍E�P������U��  ��U����ĉ�U��P�U�P�MЉH��@��������MЋU���Eԋĉ�M�P�U؉H��@����P�ݛ���E�F���E�ɉ<ȋV���U�ɉT��N���M�҉L��V���U�ɉT��EԍM�Q�N�E��-
  �U�E�P�N�U��
  �M�Q�U�R�N0�}������ ;F4u`�M��U�M�R�M���  �M�Q���  ��U���E�P�M��U��  �M�Q����  ��U��R�M��}��  �M�Q����  ����}��U�R������P�N0�}��h����;N4u`�U��E�P�M��U��_  �M�Q���  ��U���E�P�M��U��>  �M�Q���s  ��U��R�M��}��   �M�Q���U  ����U�E�P�� ���Q�N0�U������;V4�d  �E�M�Q�M��E���  �U�R���  ��M���E�Q�M��E��  �U�R����  ��M���E�Q�M��E��  �U�R��  �[����U��@���Q�M�R�U��E��E�PQR���:����M�E䍅@���P�E�Q�M�U�RPQ��������@���R�U܉E؋EP�M�QWR��������E̋F���U��M�R�������  ��U����ĉ�U��P�U�P�MЉH��@����W����MЋU���Eԋĉ�M�P�U؉H��@����P�-����M̋UЃ��E�ĉ�M؉P�U܉H��@����P�����E��F���E�ɉ<ȋV���U�ɉT��N���M�҉L��V���U�ɉT��EԍM�Q�N�E��S  �U�E�P�N�U��A  �M��U��M�R�N�/  �E�P������Q�N0�}�������;V4��   �E��M�Q�M��E���  �U�R���!  ��M���E�Q�M��E���  �U�R���   ����M��E�P�}��  �M�Q����  ��U���E�P�M��U��  �M�Q����  ����}��U�R������P�N0�}��T����;N4��   �U��E�P�M��U��G  �M�Q���|  ��U���E�P�M��U��&  �M�Q���[  ��U��R�M��}��  �M�Q���=  ��}���U�R�M��}���  �M�Q���  �����}ЋU�E�P������Q�N0�U�誢���;V4��   �E�M�Q�M��E��  �U�R����  ��M���E�Q�M��E��|  �U�R���  ��M���E�Q�M��E��[  �U�R���  ����M��E�P�}��=  �M�Q���r  ����U܍E�P������Q�N0�U������;V4��   �E؍M�Q�M��E���  �U�R���-  ��M���E�Q�M��E���  �U�R���  ��M���E�Q�M��E��  �U�R����  ����M��E�P�}��  �M�Q����  ���C;]�������@���蔓���]�����;�t!������PQ�EP������S������  �E��8�}�;���   ��    �OQ������R��莿��� ݝt����������@ݝ|����@�����P�]�Q�O����݅t����݅|����H�E��������ʋP�������H�������P�@��0����������������O�X������Q�X��݅�����X݅�����X ݅�����X(�Ⱦ���M������}�;}��4�����  �VT3�WR�ȉE��~�  ��l���蓅�����,����Pj��0�����8����e  ��;��t  ��4���� ��4����@��4����@��4����@��4����A�NH��E;���   �P��@���Q�U��@S�U�R�M��E��,���P�M�����P���{������E�PW�M�����P�M������NTPQ�9����W�M��݄��P��l�������j P��,����s���P������R��,�������W�M�跄��P��|����ۄ��j P��,����=���P��X���P��,����Z����M�"����E;FH�*���3���@��,���;�t1�F�PQ�UR���ŵ����0�����,�����,����NR�Ή�F  �M�WWW�+�  ��4����PQ�EP��,���肵����4���Q��e  �U�R�=�  �������P�}��Q�EP��������������Q��e  �� ������PQ�UR�������  �� ���P�e  �E����PQ�MQ�M��$  �U�R�{e  ��T�����;�t	P�he  ����D�����T�����X�����\���;�t	P�Ce  ���E�P��D�����H�����L����Q�EP�M��  �M�Q�e  ��_^[��]� �UR�������}�-: hH�������Pǅ����p��; �M�MQ��h���� : hH���h���Rǅh���p���: �E�MP��h�����9 hH���h���Qǅh���p��: �UR��h����}�9 hH���h���Pǅh���p��: ��U��V��FW�};�s1�;�w++���;Fu	j��������F��t*�����F_^]� ;Fu	j�������F��t���F_^]� �����������U��S�]�C�@VW��~WP������G�K�V�N�B�x u8��y u
����y t���v�N�A�x u�ȋA�x t�_�N^[]� ��v_�v^[]� ���������U��Q�UV��F�M;u;�u�������F��E�^��]� ;�t^�y ��uB�A�x u�ȋ�x u��ȋ�x t��M��A�x u;Hu�ȉM�@�x t�ER�U�R���&����M;Mu��E�^��]� ��U��Q�UV��F�M;u;�u�������F��E�^��]� ;�t^�y ��uB�A�x u�ȋ�x u��ȋ�x t��M��A�x u;Hu�ȉM�@�x t�ER�U�R��������M;Mu��E�^��]� ��U��Q�UV��F�M;u;�u���a����F��E�^��]� ;�t^�y! ��uB�A�x! u�ȋ�x! u��ȋ�x! t��M��A�x! u;Hu�ȉM�@�x! t�ER�U�R�������M;Mu��E�^��]� ��U��j�h�d�    P��SVW�`#3�P�E�d�    �e���jP�L_  �����u�3�;�t^�O��W�V�O�Nf�FH�E��UR�FP��W�������E������ƋM�d�    Y_^[��]� �M�Q��`  ��3�PP�7 �E�UR�M��
6 �E�p�hH��E�P��6 ������������U��j�h�d�    P��SVW�`#3�P�E�d�    �e���j(�|^  �����u�3�;�t^�O��W�V�O�Nf�F �E��UR�FP��W�5������E������ƋM�d�    Y_^[��]� �M�Q�`  ��3�PP�M6 �E�UR�M��:5 �E�p�hH��E�P�)6 ������������U��j�h0�d�    P��SVW�`#3�P�E�d�    �e���j�]  �����u�3�;�t^�O��W�V�O�Nf�F�E��UR�FP��W�������E������ƋM�d�    Y_^[��]� �M�Q�L_  ��3�PP�}5 �E�UR�M��j4 �E�p�hH��E�P�Y5 ������������U���SVW�}W���l�����;^t�CPW���	}����t9��W�E�M�P�ΉU��E�    �����PS�MQ��������E_^��[��]� _^�C[��]� U��j�hP�d�    P��SVW�`#3�P�E�d�    �e��ى]�C�E�}�I uO�OQ����������U�V�GH�FH�M�yI t�u��E�    V�R�������V�GP���|����F�E������E�M�d�    Y_^[��]� �M�Q�M�����j j �#4 ������U��j�hp�d�    P��SVW�`#3�P�E�d�    �e��ى]�C�E�}�! uO�OQ����������U�V�G �F �M�y! t�u��E�    V�R�������V�GP���|����F�E������E�M�d�    Y_^[��]� �M�Q�M������j j �c3 ������U��U��VW���O�A�x! ��u�
�I 9H}�@���� �x! t�;wt�;F}0�
��U��]��M�R������PV�EP���n����E_��^��]� _�F^��]� �����U��U��V��N�A�x W��u�
�I 9H}�@���� �x t�;~t�;G}2�
�U��M�R���E�    �i���PW�EP��������E_��^��]� �G_^��]� ���U��S�]�C�@VW��~WP�e����G�K�V�N�B�xI u8��yI u
����yI t���v�N�A�xI u�ȋA�xI t�_�N^[]� ��v_�v^[]� ���������U��S�]�C�@VW��~WP�����G�K�V�N�B�x! u8��y! u
����y! t���v�N�A�x! u�ȋA�x! t�_�N^[]� ��v_�v^[]� ���������U��j�h��d�    P��SVW�`#3�P�E�d�    �e���u�3��~jP��X  ��;�tf�F� �F�@�F�@�N��AH�V�BI�}��EP�������E������ƋM�d�    Y_^[��]� �M�A�PR�UR�����3�WW�0 �}�EP�M��/ �E�p�hH��M�Q�0 ���U��j�h��d�    P��SVW�`#3�P�E�d�    �e���u�3��~j(�X  ��;�tf�F� �F�@�F�@�N��A �V�B!�}��EP���@����E������ƋM�d�    Y_^[��]� �M�A�PR�UR����3�WW��/ �}�EP�M���. �E�p�hH��M�Q��/ ���U��ASVW�}=���r/�G�PQ�EP�O�:����OQ�QY  W�KY  ��h���Q- @�A�E�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z ��  �P�r;��   �v8^ u�B �F �P�R�Z �@�@�Q  ;Bu:�P�2�p�28^!u�F�p�r�q;Fu�V��p;u���V��P�P�B �P�R�Z �P�R�2�~�:�~8_!u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^ u�B �F �P�R�Z �@�@�   ;u<��r�0�r8^!u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B �P�R�Z �P�R�r�>�z�>8_!u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z �q����A�H�E�8_^�A []� ��������U��E��t�M���Q�H������]��U��QS�]�{! V�M���u=W�F�M�P������C��6PQ�MQ�K������SR��V  S��V  ���~! ��t�_^[��]� �������U���S�]�{! VW�M�t
h ��+ �M�]��ֱ����y! t�{��C�x! t���
�E�x;�ur�! �su�w�M��A9Xu�x�9u�>��~�A9u�! t���W�$����M����Q��I�M�9Yux�! t�ƉA�kW�k>  �M���A�Z�A��;Cu����! �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S �H �P �K �E��8X ��   �M��Q;z��   8_ ��   �;�ue�F�x  u�X V�F  �t����F�M��x! ut�8Z u�P8Z ta�P8Z u��Z P�@  �r>  �F�M��V �P �^ �@V�X �'����t�x  u�X V�F  �B>  ��M��x! u�P8Z u�8Z u�@  �A���v;x�J����0�8Z u�P�Z P�@  �ʱ����M��V �P �^ � V�X ��=  �_ �u��F�PQ�M�Q�N�h����VR�T  ��P�wT  �M��A��_^[��tH�A�E�M���]� �����U��Q�ыJ�A�x! S�]V��W�U��Mu-�{�} ��t9x���;x���M��t� ��@�x! t֋��}��t5�B�M;0u SVjQ���b�����E_^��@[��]� �I<  �}�U��G;C}%�MSVQ�EP���*�����E_^��@[��]� �C�PQ�UR�K�c����CP�zS  S�tS  �E���8_^�@ [��]� ���������������U��j�hФd�    P��SVW�`#3�P�E�d�    �e���j$�Q  �����u�3�;�t^�O��W�V�O�Nf�F �E��UR�FP��W�������E������ƋM�d�    Y_^[��]� �M�Q�R  ��3�PP��( �E�UR�M���' �E�p�hH��E�P��( ������������U��Q�UV��F�M;u8;�u4�@P���=����F�@�F� �F�@�N�E�F    ��^��]� ;�tb�y! ��uF�A�x! u�ȋ�x! u��I �ȋ�x! t��M��A�x! u;Hu�ȉM�@�x! t�ER�E�P�������M;Mu��E�^��]� ��U���V��~ �FW�}uW�}PjW������_^��]� S�];u&�O;K��   W�}SjW�������[��_^��]� ;�u'�@�P;W��   W�}Pj W�����[��_^��]� �G;C}M�M�]�9  �E�O9H}7�H�y! W�}��tPj W����[��_^��]� SjW�p���[��_^��]� �G9C}R�M�]�����E;Ft�O;H}7�S�z! W�}��tSj W�*���[��_^��]� PjW����[��_^��]� j W�E�P���-�����E[_�^��]� �������������U���4S�]V��W�~�G�x! u��d$ 9H}�@���� �x! t�;~t�;G��   j(�E�    �N  ������   �E� �E�@�E�@�M��A �U�B!��M�Q�MЉE������U�R���x���PW�EP��������Eԋ�}PQ�MQ�M������U�R�O  �E���PQ�EP�M��f����M�Q�}O  ���G_^[��]� �U�R�M��E�    �$ hH��E�P�E�p��% ������U��M�Ey �����%   �   @]� �   � ��������U��Vh��jah�5j�O  ������t����@ �E�F�\���^]� 3�^]� ���������������U���4Vh��jkh�5j�fO  ������t����  �ܳ�3���5�H�A�U�R�Ћ�5�Q�Jj j��E�hX�P�ы�5�B�P�M�Q�ҡ�5�H�Aj j��U�hD�R�Ћ�5�Q�J�E�P�ы�5�B�Pj j��M�h4�Q�҃�<�E�P�M���  � V�M�QPj �U�Rhy� ��� ���M�����  ��5�H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�P�M�Q�҃���^��]�����U���   ��5��P���   V�u���$hxvpi�����]ԋ�5��Q���   ���$hyvpi�����]̋�5�Q���   j hacpi���Ѓ��I  W�}���pf �����3  ��5���   �Bh�  ���Ѕ��  S���n{ Vj(���{ �?  �΋���  �M���̞��V��P����p����+  P��P���Q�U�RSV�X  ��[��~�E�P��P����1���Ou�M�薋 ��5���   ���   �Ћ�5�E����   �ȋ��   V�ЋM��Ujj QR��� �]ġ�5���   ���   �U�R������]��@q  j V�ȉE��q  �E̋}j ���\$���E��$h �  �� �M�Q�U�R�E�P���� ����   ��    �E��E��U���������Au���U�����MċM���$QV�M�譡���Mj jV�q  ��5�BH���   jV��j h  � �  ���U�R�E�P�M�Q��蚄 ��t���辄 �u��u����y j ���6z ����y j �x�  �UR�_p  ���M��E    �}� ��P��������E�PQ�EP�M������M�Q��J  ��_�   ^��]� ������U��V���= �Et	V�J  ����^]� ���������������U�조5��V��H�A�U�R�Ћ�5�Q�Jj j��E�h��P�у�j �U�Rj jj8j ���# ��5�H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�Pj j��M�h��Q�҃�j �E�Pj jj8j ���� ��5�Q�J�E�P�у�jj��� ��5�B�P�M�Q�ҡ�5�Hj j�h���A�U�R�Ѓ�j �M�Qj j jj ��� ��5�B�P�M�Q�҃�j jFjh�  ��� ��5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�у�j �U�Rj j jj ���> ��5�H�A�U�R�Ѓ�j jFjh�  ��� ��5�Q�J�E�P�ы�5�B�Pj j��M�h��Q�҃�j �E�Pj j j j ���� ��5�Q�J�E�P�ы�5�B�P�M�Q�ҡ�5�H�Aj j��U�h��R�Ѓ��M�QjjPj h�  ��� ��5�B�P�M�Q�҃����` ���Y �   ^��]����������������U�����5Vh���h  �j jh���j ��P�M�Q���E��  �E�    ��  ��j �� �\$�U�������\$�E��  ����E�    �\$� !�$R� �   ^��]��������̡�5�����������3�9(!�������U��E��pSVW��  ��;�u]h�5�E�3�P�}��]��� �   9�5��  h���h  �Sjh���SP�M�Q�Σ�5�}��]��(�  _^�C[��]� ��  ;�u(h !�U��M�R���E�    � _^�   [��]� =�  �m  h !�E��M�3�P�Ή]��x h�5�M�Q�Ή}��]��" �s ������_ ��;��'  ��5���   �Ph�  ���҅��  ����t Vj(���u ����  �M���H���V�M�����3�9(!�M���P�E�PQSV��  3ۃ�9�5~��$    �U�R�M�����C;�5|��k  j V�ȉE�k  � !�E���$PV�M��������5�QH���   jV�ЋM��j j j �k  ���Dt j ��  �MQ��j  ���M��E    蒕���E�PQ�U�R�M�蟓���E�P�VE  ��_^�   [��]� ����̋A������������̋I�   ;�u3�Ã�~�   �������U���Vj �EP���|��P�M�Q������^��]� ���������U��E@;Eu3�]�U��EHy�EH]��U����`#3ŉE��E��P�M�H�@V�U��M�E��   ;�u�   S3�W3�3ۉM�;�~�E��I �T��;�u��;Uu��A;�|�G��ȅ�y�N�;�u�O;�u3ɋL��M�O;�u3�_;�[u��y�F��D��^�M�3���! ��]ËM��E�3�^��! ��]����������������U����`#3ŉE��E��P�M�H�@�U��M�E��   ;�u�   �E�3Ʌ�~V�u9t��u��A;�|�^�M�3��x! ��]����������������U���0V�E$P�M�Q�|���U��R�E�P�|���E$�E���E�E,�E4�E�@�N�����@�N^��������������������D�E{��������������X���X��]������������P�P���]������������U��V�u�E$PV�|�����}< ��   �E���E�����E�����j" ����������D{�����E���E���E������E�E�E��������N�����N����������������n�F������^�^�F��F������������������! ����������D��{�����������N�^�N�^^]���^]Ë�^]���������U���X�`#3ŉE��ES�]VW�}3�j�}ĉ]��E��u��?  ��;���  �Eԉ �Eԉ@�Eԉ@�M��A�U��B��5�HH���   Vh�  S�҃��EȍE�P�M�QV��3���  ���  �E�C�]���E�;E��y  ���$    ��5�BH�M����   h�  Q�҃�9E��4  �ƙ�������%  ��]�yH���@����Mȿ   ��U�Q�U��Q�I�U�M�;�u�   ;�u�   �t��@����M�S�|��WV耾  �E������   �M�����3�;�u9ytk;�u	9qu3��^�A;�u9yu�   �K;�u9qu�   �;�A;�u9yu�   �(;�u9qu�   ��I;�u;�t;�u	;�u�   �E���5���Q\�J,P�E��E�P�у���uP�U�R�M��w��P�E�P�M������u�F�u�;u�������]�}ċEԋ0;�t^��$    �NQ����  �~ uA�F�x u����x u.����x t��"�F�x u��$    ;pu���@�x t���;u�u��U�R�E�PS�����  ��������EԋPQ�M�Q�M������U�R�5?  �M���_^3�[�
 ��]ÍE�P�M��u��K hH��M�Q�E�p��: �������������U���d�`#3ŉE��E�U�MS�]V�uW�}V�E��E �U��U$SV�u܉M��E��U��e�����4]���E��E� �M�WSV�b�  �E؃���2  �M���<�WSV�]������U����؋BSV�M��E��\���M��EЋA�p�~ �E�u-��    �UЋM�R�FP�P\����t�v��u�6�~ t܋E�u��E�;Ft�MЃ�PQ���\����u�E��	�V�UčEċM�9up�G��E��G��E��U�E�}��   ;�u�   3���~��$    �U�9T��u�E�@;�|�E؋M��UԉE��E��M��M�P�U��q/  �}؋u�������}� t�MԋE܋U�Q�M�PRP��c�����\���M�_^3�[�, ��]����U���  �`#3ŉE��E�M�US�]VW3�j$��t�����D����M���X�����������:  ��;���#  ������� �������@�������@�������@ �������A!j$������:  ��;���#  �� ���� �� ����@�� ����@�� ����B �� ���������@!�`Z�����`����Pj,��d�����l����R:  ��;��p#  ��h���� ��h����@��h����@��h����@(��h����A)�������Y����������@j��������������9  ��;���"  ������� �������@�������@�������A�������Bj�������9  ��;���"  ������� �������@�������@�������@�������A������VY����������@j�������������H9  ��;��f"  ������� �������@�������@�������A�������Bj�������9  ��;���!  ������� �������@�������@�������@�������A��5�BH���   Vh�  S�ы�5���BH���   Vh�  S��0����у��ˉ������a�  �ˉE��u��u��u���  ��h���;��)  �������PQ�U�R����������������P�;:  ���������PQ�M�Q������蟉��������R�:  ���������PQ�E�P�������׈��������Q��9  ���������PQ�U�R�������O���������P��9  ��h������PQ�M�Q��`����(  ��h���R�9  �� ������PQ�E�P�������_4  �� ���Q�s9  �U؋��������PQR�������74  ������P�K9  �M���_^3�[�  ��]Í������L�  ��5�QH���   h�  S�Ћ�5�QH��VP���   Wh�  S�Ѓ�P�������9�  ��D���������QSW�������������R������PV�ω�\����V�  ���p  ��������\�����T���;������*  ��T����Ǚ���4����  ��u�yO���G��5�QH���   h�  S�Ѓ�;���   ��0�������H�M��H�@�U�M�E��   ;�u�   ;�u�   W�U�R�������3  ���;l���G����t��Eԍ������uԋ|��WP��8����t3  ������V��8���Q�������Z3  ������WV�������U��j P�������H���P������R�������e�����t�����T���@��T���;������������\���������P������Q��D���R���  �������S��������a��3���$�����(�����,������������T���;��G  ���    ��T����p��P�������u��'  ��h���j�V�J  �����0����E����L0�|0Ƌ0�@�   �u�}��M�E��U�;�u�   �U��u܉}��M�E��E�    ���  �]��u��{��ǅ�y�E�HP�������nj��S�������E��_j���EӋǉEԅ�y�M�I�MԋE��\��U�@�]��E�;�u3��L��ǉM���y�B��}� �T�싽�����[�Ǎ�ݝ|����I�@���]��U��@�R�]��ݝt����Aݝ|����A��ݝ�����ݝP����AݝX����Aݝ`���u
�}� �*  ���P����D������H��H���݅D����P��L����H��P����P��0�����T���݅L����M��X��X���݅T���S�X���X�X �X(�����}� ��  �}� ��  ݅|���������������E��X�E��X�a���}� ���E��t����   �}��U���x�����x���;�si��;�wc�M�+����E�;�uF��+���=���?��  +�@��;�v*�������?+�;�s3���;�s��Q�M�������}��U���t`�Mԋ���V�M�;�uC��+���=���?�>  +�@��;�v'�������?+�;�s3���;�s��Q�M�螛���}���t��x�������}�݅P���j݅|���������Ƀ������ݕ4���݅X����E������U�݅`����E�����ݕl���݅t�������ݕH���݅|�������ݕ����݅��������ݕ���������X���X��Q����X�X����݅H�����8݅����j݅�����݅4������E���݅l�����t���������X���X��R��X�X�>�����t�����x����� �ĉ��|����P�������H�������P�H������������P��������ĉ�� ����P��$����H��(����P��,����H�P��\���P����݅|�����E��P�E�������ʋH������P������H������P�����������M��X�� ���V�X݅����X݅����X ݅����X(�����M��E�������������R��$�����������������#  �E�P�������-  ���������n  �M�SQS��`����@X�����YP��;���   ݅|���������������E��X�E��X�]^���Ű�WSRS��`�����W�����2P��݅4���ݕ,����E�ݕ4���݅l���ݕ<�������������������� ��������������Dz�������$������݅,�����݅4�����݅<�����������݅|����M��E���0�E�����W��X�X���X���X �X(�·���E�SPS��`����=W�����VO��;���   ݅|���������������E��X�E��X�Z]���M���WSQS��`�����V�����/O��݅H���ݕ���݅����ݕ���݅���ݕ�������������������� ��������������Dz�������$������݅�����݅�����݅�����������݅|����M��E���0�E�����W��X�X���X���X �X(�Ȇ���U�SRS��`����7V�����PN�����E�SPS��`����V�����6N�����̉�q�y�Y�������\����X���P���ͭ���M�SQS��`�����U������M��P������V�������U�SRS��`����U������M��P�������  ��  �M��U��<�W�ȉ�������  �������t���P��  ��5�Q\������J,WP�ыU�����S�R@S��`����E��@U�����YM��;���  ݅|���������������E��X�E��X�][���}� ���E��D�܉�8�����x����8��   �U��E��}�;�sk��;�we�Mċ�+���;�uF��+���=���?�;  +�@��;�v*�������?+�;�s3���;�s��Q�M�蛕���u��U���t�����8����S�M�;�uC��+���=���?��  +�@��;�v'�������?+�;�s3���;�s��Q�M��=����u���t�E�����u�݅t����}� ݅|�������݅|������E�R���݅�������E�����݅P�������ݕ4���݅X��������U�݅`�������ݕl���������X���X����X�X�����P�C���݅|����� ����E��E������������ʉ������,������� �������������$����X�������(����X�����݅����M��X�����݅���W�X ݅����X(范���u�WSVS��`�����R�����3K���M�Q�������(  ���=�����uJVS�������J��j P�����������P�����R����������jSVS��`����R�����K���  ��0���P��$���Q������R�U�������P��`���QVSR������ �  �E�SPS��`����HR�����aJ���}� ���E��D�܉�x����8��   �U��M��}�;�so��;�wi�M�+�����8���;�uL��+���=���?�q  +�@��;�v*�������?+�;�s3���;�s��Q�M��ђ���u��U���8�����tZ����S�M�;�uC��+���=���?�  +�@��;�v'�������?+�;�s3���;�s��Q�M��s����u���t�U�����u�݅t����}� ݅|������������݅|������E�Q���݅�������E�����݅P�������ݕ4���݅X��������U�݅`�������ݕl���������X���X��R��X�X�y��������������u��� �ĉ�� ����P��$����H��(����P��,����H�PW������P�������P���̉�P�Q�P �Q�P$�Q�P(�@,�Q�A��\���Q�Y���݅|����E��E���ʋH������P������H������P�@���� �����������������XW���X݅����X݅����X ݅����X(�V����M��U���x����������������������������R��$����$  �E�P��������$  �����������  �}�SWS��`����tO�����G��;���   ݅|���������������E��X�E��X�U����VSWS��`����0O�����iG��݅4���ݕ�����E�ݕ����݅l���ݕ���������������������C ��������������Dz�������$������݅������݅������݅������������݅|����M��E���0�E�����V��X�X���X���X �X(����u�SVS��`����tN�����F���M�SQS��`������ZN�����sF�����̉�y�Y�Y��������T����X���P���
����U�SRS��`����N�����2F��P���J���SVS��`�����M�����F��P���-��������P���  ǅ���    ��  �}� ��  ��  �MԋU��<�W�ȉ�\�����  ��\�����t���P��  ��5�Q\��\����J,WP�ыŨ�S��R�S��`���G�kM�����E��;���  ݅|���������������E��X�E��X�S����h������E��D�܉�x����0�E�j�P��8����:  �����   �U��u��u��M�;�si��;�wc�M�+����E�;�uI��+���=���?�R  +�@��;�v*�������?+�;�s3���;�s��Q�M�貍���u��U��Eԅ�tZ����S�M�;�uC��+���=���?��  +�@��;�v'�������?+�;�s3���;�s��Q�M��W����u���t�U�����u�݅P�����݅|���������݅X���Q�E������݅`������E��������݅t�������ݕH���݅|�������ݕ����݅��������ݕ���������X���X��R��X�X�\��������݅|���������� �ĉ�� ����P��$����H��(����P��,����H�P������������E��X�E��X�~����0����   󥋵8����M�V�{���E�VSPS��`����K�����XC���M�Q�������9   ���b�����uM�u�VS��$����B��j P������� ���P������R�������=���jSVS��`����J�����6C����  ��0���P��$���Q������R�U̍�����P�E���`���QRSP� ����� �  �M�SQS��`����gJ�����B��݅P���݅|�������E�݅X����D���E���x�����0݅`������E�������݅t���P����̋ă�ݕH��������݅|����u�����ݕ����݅��������ݕ���������X���X��Q��X�X�s��������������� �ĉ�� ����H��$����P��(����H��,����PV�������H�M�R�z���P���̉�P�Q�P �Q�P$�Q�P(�@,�Q�A��\���Q�U���݅|�������̉�P�Q�P�Q�P�Q�P�@�Q�A������������E��X�E��X��{����0����   �M�Q�M��`y���E��U���x�����L�����H������H���P��$�����P����.  �M�Q��������  �����������  �}�SWS��`����~H�����@��;���   ݅|���������������E��X�E��X�N��PS��RS��`����E��7H�����p@��݅H���ݝ��������݅����Pݝ �����\���݅���Qݝ(�����Z���݅|������̉�P�Q�P�Q�P�Q�P�@�Q�A������������E��X�E��X�~z����0����   �M�Q�M��x���}��U�SRS��`����G�����?��SWS��`������iG�����?�����̉�A�q�q��������M����X���P������SWS��`����+G�����D?��P���\����E�SPS��`����G�����$?��P���<�����\���Q��  ǅ\���    ���E؉E�;E�������}� �  �   �E�    �U��|��;u�u3��\��F�P�������;T������   �u�;u�u�E�    WSW��`����vF�����>��SSW��`����E��^F�����w>���MԋT�܋M��|܃��̉�Q�U؉y�Q��������L����j �M؍�   Q�������E��^W��P������R������苏����X���S违����;u�u3��D�܋�X���P������W���ܜ���E�F�N�;M�������������PQ��@���R�������n��������P�#  ��T������y! uA�A�x! u�ȋ�x! u(��ȋ�x! t���A�x! u;Hu�ȋ@�x! t��ȉ�T���;������������t����������vI���M���  �}�+}�3�����t�M����M�R�p�  F;�r싍(�����$���+θ���*���������t��S����  ��Ou�������E�;�t*��D�����    �@P����  �M��b���E�;�����u��5�QH���   j h�  S�Љ�0����������8���}�;��	  �w�ƙ�������%  �yH���@���0����+�U�Q�U��Q�I���   �U�M�;�u�   �\��@;�u3��t��G%  ���D���yH���@%  �yH���@u��D������D���WQVS��`����C������;����D���jRVS��`����C�����<��VS�������\;��j P������较��P������P�������ۍ���M��a���}�;�����������B  ��t���j Q�ȉ�<����B  �������:����4����#;����������E�;���  �P�������@�������������:�����������:����VW��`�����B�����4����P��8����H��<����P��@����@W��4�����D����:��V��4������:��W��4����E���:����tKV��4�����:����u;��<����U���t���QSRWP�54����SW�������:���H�Q��X���R����V��4����:����tNW��4����w:����u>��<����M���t���PQSVR��3���E���PV�������9���H�Q��X���R赘��V��4����):������   W��4����:�����q   ��<�����t���PSVWQ�w3����<����E���t���RPVSQ�^3����(SW��$����>9���P� ��X���RP���:����M�QV������9���P� RP�������M��t_���E�;�����������<���3�VVV�@  ��<���Q��?  ��$�������<���;�t	P�  ��������;�t	P�m  ��������������������������;�t	P�H  ���������������������������X�  �E�;�t	P�  ���������PQ��@���R�������<���������P��  ���������PQ��@���Q�������Qi��������R��  ���������PQ��@���P�������h��������Q�  ���������PQ��@���R��������h��������P�o  ��h������PQ��@���Q��`����0  ��h���R�D  �� ������PQ��@���P�������  �� ���Q�  ��@�������hx��� �M�Q��H����u��+� hH���H���RǅH���p��� �E�P��H����u���� hH���H���QǅH���p���� �U�R��H����u���� hH���H���PǅH���p��� �������������U�조5�UVj ��HH���   h�  R�ЋN����wk�$��� ��Vɉ�^]� ��VɉT�^]� �ɋT�;T�u�V�T���VɉT�^]� �ɋT�;T�u�V�T���VɉT�^]� 3� B� R� w� ����U��E��y u������y t�]�����U��E�H�y! u����H�y! t�]���̋���y! t�I�Ë�z! u�J�y! u0�ыJ�y! t��ËQ�z! u�;
u��R�z! t��y! u��������������U��M��3���tD��UUUw�I��P��  ����u(�MQ�M��E    �� hH��U�R�E�p��
� ��]� �������U��U�V�p�2�p�~! u�V�r�p�I^;Qu�A�P�B]� �J;Qu�A�P�B]� ��P�B]� ���������U��E��t�M���Q�P�I�H]��U��E��t�M��]��������������U���S�]�{) VW�M�t
h ��a� �M�]��F6����y) t�{��C�x) t���
�E�x;�ur�) �su�w�M��A9Xu�x�9u�>��~�A9u�) t���W�5���M����Q��I�M�9Yux�) t�ƉA�kW�4���M���A�Z�A��;Cu����) �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S(�H(�P(�K(�E��8X(��   �M��Q;z��   8_(��   �;�ue�F�x( u�X(V�F( �T4���F�M��x) ut�8Z(u�P8Z(ta�P8Z(u��Z(P�@( �4���F�M��V(�P(�^(�@V�X(�4���t�x( u�X(V�F( �R4����M��x) u�P8Z(u�8Z(u�@( �A���v;x�J����0�8Z(u�P�Z(P�@( �3����M��V(�P(�^(� V�X(��3���_(�M�Q��  �M��A��_^[��tH�A�E�U���]� ���U��SVW�}�) �ً�u�FP��������6W�  ���~) ��t�_^[]� ��������U��j�h�d�    PQSVW�`#3�P�E�d�    �e��E�    �]�}�u��$    ;utVWS����������}���u���E������ǋM�d�    Y_^[��]�j j �K� ��������������SVW���G�X�{ ��u�NQ���B`���6S��  ���~ ��t�G�@�G� �G�@�G    _^[����U��j�h�d�    P��SVW�`#3�P�E�d�    �e��ى]�C�E�}� uO�OQ���&J�����U�V�G�F�M�y t�u��E�    V�R�������V�GP���|����F�E������E�M�d�    Y_^[��]� �M�Q�M��__��j j �3� ������SVW���G�X�{) ��u�NQ�������6S��  ���~) ��t�G�@�G� �G�@�G    _^[����U��S�]�C�@VW��~WP������G�K�V�N�B�x u8��y u
����y t���v�N�A�x u�ȋA�x t�_�N^[]� ��v_�v^[]� ���������U��Q�UV��F�M;u;�u�������F��E�^��]� ;�t^�y) ��uB�A�x) u�ȋ�x) u��ȋ�x) t��M��A�x) u;Hu�ȉM�@�x) t�ER�U�R���v����M;Mu��E�^��]� ��U��E�UP�Ej ��Q�MQRP�������]� �����������U��j�h0�d�    P��SVW�`#3�P�E�d�    �e���}��UUUv
hx��!� �N+����*���������;�sgW�N������E��E�    P�NQ�R���S����E�������N+˸���*�����������t	S�  ���E�@�E���V����V��M�d�    Y_^[��]� �E�P�q  ��j j �� �����U��j�hP�d�    P��SVW�`#3�P�E�d�    �e���u�3��~j�$  ��;�tf�F� �F�@�F�@�N��A�V�B�}��EP���P����E������ƋM�d�    Y_^[��]� �M�A�PR�UR�]��3�WW��� �}�EP�M���� �E�p�hH��M�Q��� ���U��QVW�9+׸���*��E�������UUU+�;�s
hx��o� �Q�+׸���*���������;�v!����UUU+�;�s3���;�s��P�����_^]� ����������U��V�uW���O;�sO�;�wI+𸫪�*���������;Ou	j���I�����v���G��t?���Q�P�I�H�G_^]� ;Ou	j�������G��t���N�H�V�P�G_^]� �U��E��t�M���Q�H�����]��U��ASVW�}=���r/�G�PQ�EP�O�\���OQ�1  W�+  ��h���1� @�A�E�G�Q2�;�u�z�Q�:�A�x� 8]t�8�Q;u�:��x�Q;Bu�z�W��8Z ��  �P�r;��   �v8^ u�B �F �P�R�Z �@�@�Q  ;Bu:�P�2�p�28^!u�F�p�r�q;Fu�V��p;u���V��P�P�B �P�R�Z �P�R�2�~�:�~8_!u�W�z�~�y;Wu�w�V��   �z;Wu�w�V�   �7�V�   �68^ u�B �F �P�R�Z �@�@�   ;u<��r�0�r8^!u�F�p�r�q;Fu�V��p;Fu�V���B�P�P�B �P�R�Z �P�R�r�>�z�>8_!u�W�z�~�y;Wu�w��z;u�7��w��}�r�P8Z �q����A�H�E�8_^�A []� ��������U��j�hp�d�    P��SVW�`#3�P�E�d�    �e���j$��  �����u�3�;�t^�O��W�V�O�Nf�F �E��UR�FP��W�5������E������ƋM�d�    Y_^[��]� �M�Q�
  ��3�PP�� �E�UR�M��� �E�p�hH��E�P�� ������������U���S�]�{! VW�M�t
h ��� �M�]��fe����y! t�{��C�x! t���
�E�x;�ur�! �su�w�M��A9Xu�x�9u�>��~�A9u�! t���W�c���M����Q��I�M�9Yux�! t�ƉA�kW������M���A�Z�A��;Cu����! �pu�w�>�K�H�S�B�M��I9Yu�A��K9u���A�S�P�S �H �P �K �E��8X ��   �M��Q;z��   8_ ��   �;�ue�F�x  u�X V�F  �f���F�M��x! ut�8Z u�P8Z ta�P8Z u��Z P�@  �����F�M��V �P �^ �@V�X �e���t�x  u�X V�F  �������M��x! u�P8Z u�8Z u�@  �A���v;x�J����0�8Z u�P�Z P�@  �Ze����M��V �P �^ � V�X �q����_ �u��F�PQ�M�Q�N��V���VR�  ��P�  �M��A��_^[��tH�A�E�M���]� �����U��QS�]�{! V�M���u=W�F�M�P������C��6PQ�MQ�K�V���SR�  S�  ���~! ��t�_^[��]� �������U���V��~ �FW�}uW�}PjW�������_^��]� S�];u&�O;K��   W�}SjW�������[��_^��]� ;�u'�@�P;W��   W�}Pj W����[��_^��]� �G;C}M�M�]�g����E�O9H}7�H�y! W�}��tPj W�d���[��_^��]� SjW�P���[��_^��]� �G9C}R�M�]��a���E;Ft�O;H}7�S�z! W�}��tSj W�
���[��_^��]� PjW�����[��_^��]� j W�E�P���   ��E[_�^��]� �������������U��Q�ыJ�A�x! S�]V��W�U��Mu-�{�} ��t9x���;x���M��t� ��@�x! t֋��}��t5�B�M;0u SVjQ���R�����E_^��@[��]� �����}�U��G;C}%�MSVQ�EP��������E_^��@[��]� �C�PQ�UR�K�3T���CP�J  S�D  �E���8_^�@ [��]� ���������������U��Q�UV��F�M;u8;�u4�@P�������F�@�F� �F�@�N�E�F    ��^��]� ;�tb�y! ��uF�A�x! u�ȋ�x! u��I �ȋ�x! t��M��A�x! u;Hu�ȉM�@�x! t�ER�E�P���&����M;Mu��E�^��]� ��U���4S�]V��W�~�G�x! u��d$ 9H}�@���� �x! t�;~t�;G��   j�E�    �  ������   �E� �E�@�E�@�M��A�U�B��M�Q�MЉE��s����U�R������PW�EP���;����Eԋ�}PQ�MQ�M��R���U�R�  �E���PQ�EP�M��fR���M�Q�}  ���G_^[��]� �U�R�M��E�    �� hH��E�P�E�p��� ������U��V�u���t��5�QP��Ѓ��    ^]���������̡�5�H��@  hﾭ���Y����������U��E��t��5�QP��@  �Ѓ�]����������������U�조5�H���  ]��������������U�조5�H��  ]�������������̡�5�H��   ��U��E��t�x��u�   ]�3�]������U���s�   VW�xW�/� ������u_^]Ã} tWj V�� ��_������F��5   ^]���U���5�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�� ������u_^]�Wj V�6� ��_������F��5   ^]�������������U���5�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�3� ������u_^]�Wj V�� ��_������F��5   ^]�������������U���5�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�� ������u_^]�Wj V�6� ��_������F��5   ^]�������������U���5�E��t��s�   �I���   j j P�҃�]Ã�s�   VW�xW�3� ������u_^]�Wj V�� ��_������F��5   ^]�������������U��M��t-�=�5 t�y���A�uP��� ��]á�5�P�Q�Ѓ�]��������U��M��t-�=�5 t�y���A�uP�� ��]á�5�P�Q�Ѓ�]��������U�조5�H�U�R�Ѓ�]���������U�조5�H�U�R�Ѓ�]���������U���5�E��t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��� ������u_^]�Wj V�r� ��_������F��5   ^]���������U���5�E��tL�} t#��s�   �U�IR�URP���   �Ѓ�]Ã�s�   �U�IR�URP���  �Ѓ�]Ã�s�   VW�xW�F� ������u_^]Ã} tWj V��� ��_������F��5   ^]����������U��E��u�   ��5��t�U�IR�URP���   �Ѓ�]Ã�s�   VW�xW��� ������u_^]�Wj V�C� ��_������F��5   ^]����������U��E��u�   ��5��t,�} �U�IR�URPt���   �Ѓ�]Ë��  �Ѓ�]Ã�s�   VW�xW�-� ������u_^]�Wj V�� ��_������F��5   ^]�������U�조5�H�U�R�Ѓ�]���������U�조5�H�U�R�Ѓ�]���������U�조5�H�U�R�Ѓ�]���������U�조5�H�U�R�Ѓ�]���������U�조5�Hp�]�ࡰ5�Hp�h   �҃�������������U��V�u���t��5�QpP�B�Ѓ��    ^]���������U�조5�Pp�EP�EPQ�J�у�]� U�조5�Pp�EP�EPQ�J�у�]� U�조5�Pp�EP�EPQ�J�у�]� U�조5�Pp�EPQ�J�у�]� ��������P�P��P(�P �P�P@�P8�P0�PX�PP�PH����������X�X�����������X�X �X(���������X0�X8�X@���XH���XP�XX��������U��M�A8��   �IXV�AP�I@���I�AP�I(�AX�I ���I0���A@�I �A8�I(���IH������������Dz�u�؋��3�����^��]���W���A�IX�AP�I�A8�I�A�I@�AP�I@�U��A8�IX�]������IH�����I0�����e��	����ݝx����A�I(�U��A�I �U��AX�I �]��AP�I(�����IH�E����	���������I�������]��A8�I(�A@�I �����	�������I���E��e��I0�������]��E��e����]����e��ˋE��x������]������]��AH�I@�A0�IX�����]��AX�I�AH�I(�����]��A0�I(�A@�I�����]��AP�I0�AH�I8�����]��AH�I �AP�I�����]��A8�I�A0�I �   �����]��_^��]�����U��y0 ts��U�����Au���A�Z����Au�B�Y�A�Z����Au�B�Y�A�����z��Y�A �Z����z�B�Y �A(�Z����zZ�B�Y(]� �E��Q�P�Q�P�Q �P�Q$�P�Q(�@�A,�Q�A��Q �A�A$�Q�Q(�A�A,�Q�A�A0   ]� ��3ɉ�H�H�H�V��V�7����FP�.���3����F�F^��3���A�A�A����A�`�
�@�b�	���B�a�������U����   ��UV���q�U�W3��<��M��}��'	  S�]����  ��؋���M�U��>���U�@�U���� �U��@�@�B�@�������@���@�   ���]��E��U�;���  �w�����  �w�������F�܍B��   �U������������ˋP��R�э����]��B���B�P���R���U����E������]��E��M��E������������]��E����E����E��E��]����E��]����E��]����]����U��E��U�����B���B���U������������]��E����E����������E������E��E��]����E��]����E��]��]��U���E��U��R�э����N�B���B�P���R���U������������]��E����E����������E������E��E��]����E��]����E��]����U��E��]�����B���B���U����E��������]��E����E����������E������E��E��U����E��]����E��U��E��U��T����E�ɋU�����������;���   �ߍ���+�������͋�@�������O�]��@���]��@���U������M������]��E��E����E������E����������E��E��U����E��]����E��U��E��E��U�u�������������������������[�[�E������������������ ��������������Dz���������E��+������������������M����M��E������������������[H���[P���[X�E����E���������zu������������zh�����CP���CX���CH���CX�������cH���[���[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@��   ������������z]�CX���CP�����cH�CH���CP�������[�[ �[(�C(�KP�C �KX���CX�K�C(�KH���CH�K �CP�K�����[0�[8�[@�]�CP���CX�����CH���CX�����cP���[0���[8�[@�C8�KX�C@�KP���CH�K@�C0�KX���C0�KP�C8�KH�����[�[ �[(��$���SQ�����E��U�   �����}��M������3�3��u��u���|)�A�����B�4�u�0u��u�p��J�u�u�U�E;�}�Q���E���u��U��1���@���K�I�E    ��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�@�K@���CX�H�D��@�����U���]�� �K��C0�H���@�KH��� �K �C�@�K8���@�KP��� �K(�C�C@�H���CX�H���U����n  �A�������@�E����E   �E�
���������ɋEH���׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E������������������������������E����]��E��]����]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H�E@������]������M������������������������]��E��]��E��]�׋��@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������]��E�E����]���E����]��E��M����@�E�Ѝ��K��C0�H���CH�H��� �K �C�@�K8���@�KP���C(��C�C@�H���CX�H���]������M������������������������U��E��]��E��U������������������9M|��[��_��^���؋�]� ���������ʋE�����׋��@�E�Ѝ��K��C0�H���CH�H���]�� �K �C�@�K8���@�KP���]��C(��C�C@�H���CX�H�E@�E���]����E��������������������M����������]��E��E�;��T�����[������_��^��]� �����h�5Ph_� �@0 ���������������h�5jh_� �0 ����uË@����U��V�u�> t/h�5jh_� ��/ ����t��U�M�@R�Ѓ��    ^]���U��Vh�5jh_� ���/ ����t�@��t�MQ����^]� 3�^]� �������U��Vh�5jh_� ���y/ ����t�@��t�MQ����^]� 3�^]� �������U��Vh�5jh_� ���9/ ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5jh_� ����. ����t�@��t�MQ����^]� 3�^]� �������U��Vh�5j h_� ���. ����t�@ ��t�MQ����^]� 3�^]� �������U��Vh�5j$h_� ���i. ����t�@$��t�MQ����^]� 2�^]� �������Vh�5j(h_� ���,. ����t�@(��t��^��3�^������Vh�5j,h_� ����- ����t�@,��t��^��3�^������U��Vh�5j0h_� ����- ����t�@0��t�MQ����^]� 3�^]� �������U��Vh�5j4h_� ���- ����t�@4��t�M�UQR����^]� ���^]� ��Vh�5j8h_� ���L- ����t�@8��t��^��3�^������U��Vh�5j<h_� ���- ����t�@<��t�MQ����^]� ��������������U��Vh�5j@h_� ����, ����t�@@��t�MQ����^]� ��������������U��Vh�5jDh_� ���, ����t�@D��t�MQ����^]� 3�^]� �������U��Vh�5jHh_� ���Y, ����t�@H��t�MQ����^]� ��������������Vh�5jLh_� ���, ����t�@L��t��^��3�^������Vh�5jPh_� ����+ ����t�@P��t��^��3�^������Vh�5jTh_� ���+ ����t�@T��t��^��^��������Vh�5jXh_� ���+ ����t�@X��t��^��^��������Vh�5j\h_� ���\+ ����t�@\��t��^��^��������U��Vh�5j`h_� ���)+ ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�5jdh_� ����* ����t�@d��t�M�UQR����^]� 3�^]� ���U��Vh�5jhh_� ���* ����t�@h��t�M�UQ�MR�UQ�MRQ����^]� ��������������U��Vh�5jlh_� ���Y* ����t�@l��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5jph_� ���	* ����t�@p��t�M�UQR����^]� 3�^]� ���U��Vh�5jth_� ����) ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�5jxh_� ���) ����t�@x��t�M�UQR����^]� 3�^]� ���U��Vh�5j|h_� ���I) ����t�@|��t�MQ����^]� 3�^]� �������U��Vh�5h�   h_� ���) ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h_� ���( ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�5h�   h_� ���V( ����t+���   ��t!�M�UQ�MR�UQ�MR�UQR����^]� ���^]� ������������U��Vh�5h�   h_� ����' ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U���|��A���U����U����U���  S�V�E��EW�����������   ���������U�r�z�
�R;��4v���4��I�$ȍ��F�R�a���F�a�uB�!�]��B�a�U��B�a�U������������]��E����E����������E��������E��G��$ȍ��]��B�a�U��B�a�U������������]��E����E����������E��������E��������M�������_�U�^��[�U����U��������������������� ��������������D�Ez���P�P���]� �������E�����E����X�M��X��]� ����U���@����A���E�    �����]����]��]�����������]����]��]����   �	S�]VW�M��E����������t[��%�����E�M�����@��P������F�@��R�M������~���Q�M������v;�t�v��P�M������M����M��M�u��}� _^[tV�E؋E�E����E��E����E��E����@�������������X���X��� ���`���`�E����X�X��]� ��E����������P���P�E����X�X��]� �����������̋Q3���|�	��t��~�    t@��Ju��3�����������U��QV�u��;�}�	���    u@��;�|����^]� +�@^]� �����������U��VW�}��x+�1��t%�Q3���~�΍I �1�������;�t@��;�|���_^]� �Q3���~!V�1�d$ ���   @u	�����t@��Ju�^�����̋QV3���~�	�d$ ����ШtF��Ju��^�����������U��Q3�9A~��I ��$������@;A|�Q��~YSVW�   3ۋ���x5��%����E���;�}$�I �������%���;E�u�
   �F;q|ߋQG�G���;�|�_^[��]�����������U��	����%�����E��   @t������A��wg�$�X�E�M� �������]� ��M��P�E�]� �H�U�
�@�M�]� �P�M��P�E�]� �H�U�
� �M�]� ���/C����U����S��V�����W�   @t���������];�t�����u�};�tK�����tC��}�����t�������t�Ӄ��t��_%   ��^�[]� �%   ���   @�_^[]� ����V��V�'����FP����3����F�F^��U��SV��WV�����^S������E3����~�~;�t_��5�Q���   h����jIP�у��;�t9�}��t;��5�B���   h����    jNQ�҃����uV������_^3�[]� �E�~_�F^�   []� ����������U��V��WV�S����FP�J����}���F    �F    ����   �? ��   �G����   ��5�Q���  h����jlP�у����t>� t@�G��t9��5�Jh����    ���  jqR�Ѓ��F��u���v���_3�^]� �O��N�G�F��    ���t��t��tQPR�� ���F��t�VP��RP�GP�  ��_�   ^]� ��������U��SV��WV�B����~W�9���3����F�F9E�  �];���   ��5�Qh����    h�   P���  �Ѓ����t@�} tN�]��tD��5�Q���  h����    h�   P�у����u���n���_^3�[]� �^�]�0�]�F   ��5�B���  h��h�   j�у����t���^��t��    ��t�UQRP��� ���E��t!�N�?�W�QWP�R  ��_^�   []� ��_^�   []� ���U��Q�A�E� ��~JS�]V�1W����$    ����������;�u�   @u�����u3��	�   ����U���Ou�_^[�E��Ћ�]� �����������U��S�]V��3�W�~���F�F�CV;C��   �t���W�n���3��F�F��5�Q���   h��jIj�Ѓ������   ��5�Q���   h��jNj�Ѓ����uV������_��^[]� ��F   �F   ����K�H�C��B�_��^�   []� �����W�����3��F�F��5�B���   h��jIj�у����t[��5�B���   h��jNj�у�����\�����F   �F   ����S�Q��K�H��C�B��   _��^[]� �����������U��3�V���F�F�F�EP������^]� �������������U��EVP��������^]� ����������U��U��t�M��t�E��tPRQ�P� ��]������������h�5Ph� �` ���������������h�5jh� �? ����uË@����U��V�u�> t/h�5jh� � ����t��U�M�@R�Ѓ��    ^]���U��Vh�5jh� ���� ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh�5jh� ��� ����t�@��t�M�UQR����^]� 3�^]� ���U��Vh�5jh� ���Y ����t�@��t�M�UQ�MRQ����^]� 3�^]� ���������������Vh�5jh� ��� ����t�@��t��^��^��������U��Vh�5j h� ���� ����t�@ ��t�MQ����^]� ��������������U��Vh�5j$h� ��� ����t�@$��t�M�UQR����^]� 3�^]� ���U��Vh�5j(h� ���Y ����t�@(��t�M�UQR����^]� 3�^]� ���U��Vh�5j,h� ��� ����t�@,��t�M�UQR����^]� 3�^]� ���U��Vh�5j0h� ���� ����t�@0��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5j4h� ��� ����t �@4��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5j8h� ���9 ����t%�@8��t�M�E�UQ�M���$RQ����^]� 3�^]� ������U��Vh�5j@h� ���� ����t�@@��t�M�UQR����^]� 3�^]� ���U��Vh�5jDh� ��� ����t�@D��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5jHh� ���Y ����t �@H��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jLh� ���	 ����t�@L��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5jPh� ��� ����t�@P��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5jTh� ���i ����t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jXh� ��� ����t �@X��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jdh� ���� ����t%�@d��t�E�M�U���$Q�MRQ����^]� 3�^]� ������U��Vh�5jhh� ���y ����t �@h��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jlh� ���) ����t$�@l��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�5jph� ���� ����t �@p��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jth� ��� ����t�@t��t�M�UQR����^]� 3�^]� ���U��Vh�5jxh� ���I ����t �@x��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5j|h� ���� ����t�@|��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5h�   h� ��� ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h�   h� ���V ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h� ��� ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h� ��� ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h�   h� ���f ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h�   h� ��� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���v ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h�   h� ���& ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���6 ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h� ���F ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5j\h� ���� ����t�@\��t�M�UQ�MRQ����^]� 3�^]� ���������������U��Vh�5j`h� ��� ����t�@`��t�M�UQR����^]� 3�^]� ���U��Vh�5j<h� ���i ����t$�@<��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�5h�   h� ��� ����t���   ��t�MQ����^]� 3�^]� �U��Vh�5h�   h� ���� ����t���   ��t�MQ����^]� 3�^]� �U��Vh�5h�   h� ��� ����t'���   ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh�5h�   h� ���F ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t#���   ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h�   h� ���V ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h� ��� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ���f ����t,���   ��t"�E�M�U���$Q�MR�UQR����^]� 3�^]� ������������U��Vh�5h�   h� ��� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t���   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h�   h� ���f ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ��� ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   h� ����
 ����tG���   ��t=�E(�MP���ĉ�M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�$ 3�^]�$ �U��Vh�5h�   h� ���V
 ����tN���   ��tD�E0�E(�MP�� ���\$��M�H�M�H�M�H�M �H�M$�H�E�MPQ����^]�, 3�^]�, ����������U��Vh�5h�   h� ����	 ����t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h   h� ���	 ����t��   ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h  h� ���6	 ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h  h� ���� ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h  h� ��� ����t��  ��t�M�UQR����^]� 3�^]� �������������U��Vh�5h  h� ���F ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh�5h  h� ���� ����t#��  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h  h� ��� ����t'��  ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �U��Vh�5h  h� ���V ����t��  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h   h� ��� ����t��   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h$  h� ��� ����t#��$  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h(  h� ���f ����t#��(  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h,  h� ��� ����t3��,  ��t)�M$�U Q�MR�UQ�MR�UQ�MR�UQR����^]�  3�^]�  �����U��Vh�5h0  h� ��� ����t��0  ��t�MQ����^]� ��������U��Vh�5h4  h� ���v ����t��4  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h8  h� ���& ����t��8  ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h<  h� ���� ����t#��<  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5h@  h� ��� ����t#��@  ��t�M�UQ�MR�UQR����^]� 3�^]� �����U��Vh�5hD  h� ���6 ����t��D  ��t�M�UQ�MRQ����^]� U��Vh�5hH  h� ���� ����t��H  ��t�M�UQ�MRQ����^]� U���V��FT��u
���^��]� �V$�MjRP�E�M�P�M��E��� ��t�+FT^����]� �����U���V��FX��u
���^��]� �V(�MjRP�E�M�P�M��E��� ��t�+FX^����]� �����U���V��F\��u
���^��]� �V,�MjRP�E�M�P�M��E���f ��t�+F\^����]� �����U���V��FL��u
���^��]� �V4�MjRP�E�M�P�M��E���E������ ��t�+FL^����]� ��������������U���V��F<��u
���^��]� �V$�MjRP�E�M�P�M��E��� ��t�+F<^����]� �����U���V��F@��u
���^��]� �V(�MjRP�E�M�P�M��E���f ��t�+F@^����]� �����U���V��FD��u
���^��]� �V,�MjRP�E�M�P�M��E��� ��t�+FD^����]� �����U���V��FP��u
���^��]� �V �MjRP�E�M�P�M��E���� ��t�+FP^����]� �����U���V��FH��u
���^��]� �V0�MjRP�E�M�P�M��E���E������o ��t�+FH^����]� ��������������U���V��F8��u
���^��]� �V �MjRP�E�M�P�M��E��� ��t�+F8^����]� �����U��E�@�M+A]� �������������U��E��5� ]��U�조5�P8�EPQ�JD�у�]� ���̡�5�H8�Q<�����U�조5�H8�A@V�u�R�Ѓ��    ^]�������������̡�5�H8�������U�조5�H8�AV�u�R�Ѓ��    ^]��������������U�조5�P8�EP�EP�EPQ�J�у�]� ������������U�조5�P8�EP�EPQ�J�у�]� ��5�P8�BQ�Ѓ����������������U�조5�P8�EPQ�J �у�]� ����U�조5�P8�EP�EP�EP�EP�EPQ�J$�у�]� ����U�조5�P8�EP�EP�EP�EP�EP�EPQ�J�у�]� U�조5�P8�EP�EPQ�J(�у�]� U�조5�P8�EP�EP�EPQ�J,�у�]� ������������U�조5�P8�EP�EP�EPQ�J�у�]� ������������U�조5�P8�EP�EP�EP�EP�EPQ�J�у�]� ����U�조5�P8�EP�EPQ�J0�у�]� U�조5�P8�EP�EP�EPQ�J4�у�]� ������������U�조5�P8�EPQ�J8�у�]� ����U�조5�H��x  ]��������������U�조5�H��|  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H�A,]�����������������U�조5�H�QV�uV�ҡ�5�H�Q8V�҃���^]�����̡�5�H�Q<�����U�조5�H�I@]����������������̡�5�H�QD����̡�5�H�QH�����U�조5�H�AL]�����������������U�조5�H�IP]�����������������U�조5�H��<  ]��������������U�조5�H��,  ]��������������U�조5�H�E���   �PPR�P@R�P0R�P R�PRP�EP�у�]������������̡�5�H���   �⡰5�H���  ��U�조5�H�U�ER�UP�ER�UP���   Rh�.  �Ѓ�]����������������U�조5�H�A]�����������������U�조5�H��\  ]��������������U�조5�H�AT]�����������������U�조5�H�AX]�����������������U�조5�H�A\]����������������̡�5�H�Q`����̡�5�H�Qd����̡�5�H�Qh�����U�조5�H�Al]�����������������U�조5�H�Ap]�����������������U�조5�H�At]�����������������U�조5�H��D  ]��������������U�조5�H��  ]��������������U�조5�H�Ix]�����������������U�조5�H��@  ]��������������U��V�u���"  ��5�H�U�A|VR�Ѓ���^]���������U�조5�H���   ]��������������U�조5�H��h  ]��������������U�조5�H��d  ]��������������U�조5�H���  ]�������������̡�5�H���   ��U�조5�H��l  ]��������������U�조5�H��   ]��������������U�조5�H��  ]��������������U��V�u����  ��5�H���   V�҃���^]���������̡�5�H��`  ��U�조5�H��  ]��������������U�조5�H�U���   ��R�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]�����U�조5�H���  ]��������������U��U�E��5�H�E���   R���\$�E�$P�у�]�U�조5�H���   ]��������������U�조5�H���   ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���   ]��������������U�조5�H���   ]��������������U�조5�H���   ]��������������U�조5�H���   ]��������������U�조5�H���   ]��������������U�조5�H���   ]��������������U�����5�P�E�P�E�P�E�PQ���   �у����#E���]����������������U�����5�P�E�P�E�P�E�PQ���   �у����#E���]����������������U�����5�P�E�P�E�P�E�PQ���   �у����#E���]����������������U�조5�H��8  ]��������������U��V�u(V�u$�E�@��5�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U��V�u(V�u$�E�@��5�R0V�u V�uV�uV�uV�uV�uVP���   Q�Ѓ�(^]�$ �����������U�조5�P0�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���   �у�(]�$ �U�조5�P0�EP�EP�EP�EPQ���   �у�]� ����̡�5�P0���   Q�Ѓ�������������U�조5�P0�EP�EPQ���   �у�]� �������������U�조5�P0�EP�EP�EP�EPQ���   �у�]� ����̡�5�P0���   Q�Ѓ������������̡�5�H0���   ��U�조5�H0���   V�u�R�Ѓ��    ^]�����������U�조5�H��H  ]��������������U�조5�H��T  ]�������������̡�5�H��p  �⡰5�H���  ��U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H�U�E��X  ��VR�UPR�E�P�ыu�    �F    ��5���   �Qj PV�ҡ�5���   ��U�R�Ѓ� ��^��]��������U���4VhLGOg�M���  ��5�Q��X  3�VP�E�hicMCP�ы�5�u��u����   VP�A�U�R�Ћ�5���   �
�E�P�у� �M��r�  ��5���   �PT�M�Q�҃���u'�u�����  ��5���   ��U�R�Ѓ���^��]Ë�5���   �JT�E�P�ыu��P�����  ��5���   ��M�Q�҃���^��]���������������U�조5�H��  ]��������������U�조5�H��\  ]��������������U�조5�H�U��t  ��V�uVR�E�P�у�����  �M����  ��^��]�����U�조5�H�U���  ��VWR�E�P�ы�5�u���B�HV�ы�5�B�HVW�ы�5�B�P�M�Q�҃�_��^��]����������������U�조5�H�U���  ��VWR�E�P�ы�5�u���B�HV�ы�5�B�HVW�ы�5�B�P�M�Q�҃�_��^��]����������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H�U�E��VWj R�UP�ERP��t  �U�R�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�(_��^��]��U�조5�H�U�E��VR�UP�ERP���  �U�R�Ћu�    �F    ��5���   j P�BV�Ћ�5���   �
�E�P�у�$��^��]���U�조5�H��8  ]��������������U���  �`#3ŉE��M�EPQ������h   R��� ����x	=�  |#���5�H��0  h�hF  �҃��E� ��5�H��4  ������Rh`��ЋM�3̓�迉 ��]�������U�조5�H��  ��V�U�WR�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�_��^��]����U�조5�H��  ��V�U�WR�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�_��^��]����U�조5�H��p  ��4�҅���   h���M��%�  ��5�P�E�R4Ph���M��ҡ�5�P�E�R4Ph���M��ҡ�5�H��X  j �U�R�E�hicMCP�ы�5�E�    �E�    ���   j P�A�U�R�Ћ�5���   �
�E�P�ы�5���   ��M�Q�҃�$�M���  ��]��������U�조5�H��p  ��4V�҅�u��5�H�u�QV�҃���^��]�Wh!���M��,�  ��5�P�E�R4Ph!���M��ҡ�5�H��X  3�V�U�R�E�hicMCP�ы�5�u��u����   VP�A�U�R�Ћ�5���   �
�E�P�ы�5���   �PH�M�Q�ҋu����5�H�QV�ҡ�5�H�QVW�ҡ�5���   ��U�R�Ѓ�4�M���  _��^��]������U�조5�H��p  ��4V�҅�u��5�H�u�QV�҃���^��]�Wh����M���  ��5�P�E�R4Ph����M��ҡ�5�H��X  3�V�U�R�E�hicMCP�ы�5�u��u����   VP�A�U�R�Ћ�5���   �
�E�P�ы�5���   �PH�M�Q�ҋu����5�H�QV�ҡ�5�H�QVW�ҡ�5���   ��U�R�Ѓ�4�M���  _��^��]������U�조5�H��p  ��4�҅�u��]�Vh#���M��$�  ��5�P�E�R4Ph#���M��ҡ�5�H��X  3�V�U�R�E�hicMCP�ы�5�u��u����   VP�A�U�R�Ћ�5���   �
�E�P�ы�5���   �P8�M�Q�ҋ�5���   ��U�R�Ѓ�(�M����  ��^��]���������������U�조5�H��p  ��4�҅�u��]�Vhs���M��D�  ��5�P�E�R4Phs���M��ҡ�5�H��X  3�V�U�R�E�hicMCP�ы�5�u��u����   VP�A�U�R�Ћ�5���   �
�E�P�ы�5���   �P8�M�Q�ҋ�5���   ��U�R�Ѓ�(�M����  ��^��]���������������U�조5�H���  ]��������������U�조5�H��@  ]��������������U�조5�H���  ]��������������U��V�u���t��5�QP��D  �Ѓ��    ^]������U�조5�H��H  ]��������������U�조5�H��L  ]��������������U�조5�H��P  ]��������������U�조5�H��T  ]��������������U�조5�H��X  ]��������������U�조5�H��\  ]�������������̡�5�H��d  ��U�조5�H��h  ]��������������U�조5�H��l  ]�������������̡�5�H���  ��U�조5�H�U���  ��VR�E�P�ыu��P�����  �M����  ��^��]�����U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�H��$  ]��������������U�조5�H��(  ]��������������U�조5�H��,  ]�������������̡�5�H��0  �⡰5�H��<  ��U�조5�H���  ]�������������̡�5�H���  ��U�조5�H���  ]������������������������������U�조5�H��  ]�������������̡�5�H��P  �⡰5���   ���   ��Q��Y��������U�조5�H�A�U��� R�Ћ�5�Q�Jj j��E�hd�P�ы�5�B�P�M�Q�ҡ�5�H�I�U�R�E�P�ы�5�B�P<�� �M��ҋ�5�Q�M�RLj�j�QP�M��ҡ�5�H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�P�M�Q�҃���]��������������U��E��u��5�MP�EPQ�c ��]��������������̋�3ɉ�H�H�H�U��V��~ W�}u3hh�j;h�5j轡������t
W����  �3��F��u_^]� �~ t3�9_��^]� ��5�H<�W�҃�3Ʌ����_�F   ^��]� ��V���F   ��5�H<�Q��3Ʌ����^��������������̃y t�   ËA��uË�5�R<P��JP�у��������U����u��5�H�]� ��5�J<�URP�A�Ѓ�]� ���������������U�존5��u��5�H�]Ë�5�J<�URP�A�Ѓ�]�U�존5��$V��u��5�H�1���5�J<�URP�A�Ѓ�����5�Q�J�E�SP�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@�� j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у���[t.��5�B�u�HV�ы�5�B�P�M�Q�҃���^��]á�5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�u�QV�ҡ�5�H�A�U�VR�Ћ�5�Q�J�E�P�у���^��]���������������U�존5��$SV��u��5�H�1���5�J<�URP�A�Ѓ�����5�Q�J�E�P�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@�� j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у���t/��5�B�u�HV�ы�5�B�P�M�Q�҃���^[��]á�5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����3�����5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�u�QV�ҡ�5�H�A�U�VR�Ћ�5�Q�J�E�P�у���^[��]����������������U�존5��$SV��u��5�H�1���5�J<�URP�A�Ѓ�����5�Q�J�E�P�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@�� j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у���t/��5�B�u�HV�ы�5�B�P�M�Q�҃���^[��]á�5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����3�����5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����������5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�u�QV�ҡ�5�H�A�U�VR�Ћ�5�Q�J�E�P�у���^[��]��U�존5��$SV��u��5�H�1���5�J<�URP�A�Ѓ�����5�Q�J�E�P�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@�� j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у���t/��5�B�u�HV�ы�5�B�P�M�Q�҃���^[��]á�5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����3�����5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����������5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�A�U�R�Ћ�5�Q�Jj j��E�h��P�ы�5�B�@@��j �M�Q�U�R�M��Ћ�5�Q�J���E�P���у����������5�P�E��RHjP�M��ҡ�5�P�E�M��RLj�j�PQ�M��ҡ�5�H�u�QV�ҡ�5�H�A�U�VR�Ћ�5�Q�J�E�P�у���^[��]����U�조5�H<�A]����������������̡�5�H<�Q�����V��~ u>���t��5�Q<P�B�Ѓ��    W�~��t���
�  W�������F    _^��������U���V�E�P���>�  ��P�������M�����  ��^��]��̃=�5 uK��5��t��5�Q<P�B�Ѓ���5    ��5��tV����  V�z�������5    ^������������U���H��5�H�AS�U�V3�R�]��Ћ�5�Q�JSj��E�h��P�ы�5�B<�P�M�Q�ҋ�5�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]��H �M�Q�U�R�M�� ���&  W�}�}���   ��5���   �U��ATR�Ћ�������   ��5�Q�J�E�P���ы�5�B���   ���M�Qj�U�R���Ћ�5�Q�J���E�P�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Bx��W�M����E���t�E� ��t��5�Q�J�E�P����у���t��5�B�P�M�Q����҃��}� u"�E�P�M�Q�M�� ��������E�_^[��]ËU��U�_�E�^[��]��U���DSV�u3ۉ]�;�u_��5�H�A�U�R�Ћ�5�Q�JSj��E�h��P�ы�5�B<�P�M�Q�ҋ�5�H�A�U�R�Ѓ�;�u^3�[��]�V�M�]�� �M�Q�U�R�M��� ���p  W�}��I �E����   ��5���   �U��ATR�Ћ�������   ��5�Q�J�E�P���ы�5�B���   ���M�Qj�U�R���Ћ�5�Q�J���E�P�ы�5�B�P�M�QV�ҡ�5�H�A�U�R�Ћ�5�Q�Bx��W�M����E��t�E ��t��5�Q�J�E�P����у���t��5�B�P�M�Q����҃��} tC�E�_^�E�[��]Ã�u1�E���t*��5���   P�BH�Ћ�5�Q���ȋBxW�Ѕ�t"�M�Q�U�R�M��r ��������E�_^[��]ËM��M�_�E�^[��]�U��E��V3�;���   P�M��� �EP�M�Q�M�u��u� ����   �u���E���tA��t<��uZ��5���   �M�PHQ�ҋ�5�Q���ȋBxV�Ѕ�u-�   ^��]Ë�5���   �E�JTP��VP�[�������uӍUR�E�P�M�� ��u�3�^��]����������V��~ u>���t��5�Q<P�B�Ѓ��    W�~��t����  W脐�����F    _^��������U�조5�E�PH�B���$Q�Ѓ�]� ���������������U�조5�PH�EPQ���   �у�]� �U�조5�PH�EPQ���  �у�]� �U�조5�PH�EPQ���  �у�]� �U�조5�PH�EP�EPQ��  �у�]� �������������U�조5�PH�EP�EPQ��  �у�]� ������������̡�5�PH���  Q�Ѓ�������������U�조5�PH�EPQ���  �у�]� ̡�5�PH���   j Q�Ѓ�����������U�조5�PH�EPj Q���   �у�]� ��������������̡�5�PH���   jQ�Ѓ�����������U�조5�PH�EPjQ���   �у�]� ��������������̡�5�PH���   jQ�Ѓ����������U�조5�PH�EPjQ���   �у�]� ���������������U�조5�PH�EP�EPQ���   �у�]� �������������U�조5�PH�EP�EPQ���   �у�]� ������������̡�5�PH���   Q�Ѓ�������������U�조5�PH�EP�EP�EP�EP�EPQ���  �у�]� �U��EVWP����6  ������t�E��5�QH���   PVW�у���_^]� �����U��EVW���MPQ��6  ������t�M��5�BH���   QVW�҃���_^]� ̡�5�PH���   Q�Ѓ������������̡�5�PH���   Q�Ѓ�������������U�조5�PH�EPQ���   �у�]� �U�조5�PH�EPQ���   �у�]� �U�조5�PH�EP�EPQ��8  �у�]� �������������U�조5�PH�EP�EPQ��   �у�]� ������������̡�5�PH���  Q�Ѓ������������̡�5�PH���  Q�Ѓ������������̡�5�PH���  Q�Ѓ������������̡�5�PH��  Q�Ѓ������������̡�5�PH��  Q�Ѓ�������������U�조5�PH�EP�EPQ��  �у�]� �������������U�조5�PH�EP�EP�EPQ��   �у�]� ���������U�조5�PH�EP�EP�EP�EPQ��|  �у�]� �����U�조5�PH�EPQ��  �у�]� ̡�5�PH��T  Q�Ѓ�������������U�조5�PH�EP�EPQ��  �у�]� �������������U�조5�PH�EPQ��8  �у�]� �U�조5�PH�EPQ��<  �у�]� �U�조5�PH�EPQ��@  �у�]� �U�조5�PH�EP�EP�EPQ��D  �у�]� ��������̡�5�PH��L  Q��Y��������������U�조5�PH�EPQ��H  �у�]� ̡�5V��H@�Q,WV�ҋ�5�Q��j �ȋ��   h�  �Ћ�5�QH�����   h�  V�Ѓ���
��t_3�^Ë�_^�̡�5�P@�B,Q�Ћ�5�Q��j �ȋ��   h�  �������U�조5�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�조5�E�PH�E��  ��P�EP���$Q�M�Q�ҋM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����U�조5�PH�EP�EP�EPQ��   �у�]� ��������̡�5�HH��  ��U�조5�HH��  ]��������������U�조5�E�PH��$  ���$Q�Ѓ�]� �����������̡�5�PH��(  Q�Ѓ�������������U�조5�PH�EP�EPQ��,  �у�]� �������������U�조5�E�PH�EP�E���$PQ��0  �у�]� ���̡�5�PH���  Q�Ѓ������������̡�5�PH��4  Q�Ѓ������������̋��     �������̡�5�PH���|  jP�у���������U�조5�UV��HH��x  R��3Ƀ������^��]� ��̡�5�PH���|  j P�у��������̡�5�PH��P  Q�Ѓ������������̡�5�PH��T  Q�Ѓ������������̡�5�PH��X  Q�Ѓ�������������U�조5�PH��Q��\  �E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ����̡�5�PH��`  Q�Ѓ�������������U�조5�PH�EPQ��d  �у�]� �U�조5�E�PH��h  ���$Q�Ѓ�]� ������������U�조5�E�PH��t  ���$Q�Ѓ�]� ������������U�조5�E�PH��l  ���$Q�Ѓ�]� ������������U�조5�PH�EPQ��p  �у�]� �U�조5�PH�EP�EP�EP�EPQ���  �у�]� �����U�조5�PH�EP�EP�EP�EP�EP�EPQ���  �у�]� �������������U�조5�E�HH�U �ER�UP�E���$R�UP���   R�Ѓ�]������������U��U�E��5�HH�E���   R�U���$P�ERP�у�]����������������U���E�M�ȵ�,m �M;�|�M;�~��]�����������U�조5�PH�E���   Q�MPQ�҃�]� ������������̡�5�PH���   Q��Y�������������̡�5�PH���   Q�Ѓ������������̡�5�PH���   Q��Y��������������U�조5�PH�EP�EPQ���   �у�]� �������������U�조5�PH�EP�EP�EP�EP�EPQ���  �у�]� ̡�5�PH��t  Q��Y�������������̋�� Ե�@    ��Ե��5�Pl�A�JP��Y��������U�조5V��Hl�V�AR�ЋE����u
�   ^]� ��5�Ql�MQ�MQ�
P�EP��3҃����F^��]� ������̋A��uË�5�QlP�B�Ѓ�������U�조5�Pl�I�R�EP�EP�EP�EPQ�ҋE�M��;�u�E]� 9Mt���]� ������������U��U�E��5�HH�ER�U���$P���  R�Ѓ�]����U�조5�HH���  ]��������������U�조5�HH���  ]��������������U��U0�E(��5�HH�E$R�U ���$P�ER�UP�ER�UP�ER�UP���  R�Ѓ�,]������������U�조5�HH���  ]��������������U�조5�E�PH�EP���$Q���  �у�]� ��������U���SV���!  �؉]����   �} ��   ��5�HH��p  j h�  V�҃��E��u
^��[��]� �MW3��}��0  ����   �]��I �E�P�M�Q�MW��  ��t_�u�;u�W�I ������u�E����ҋL�;L�t-��5�Bl�S�@����QR�ЋD������t	�M�P��  F;u�~��}��MG�}��  ;��x����]�_^��[��]� ^3�[��]� U�����5SV�ًHH��p  j h�  S�]��ҋ�����u
^3�[��]� �E��u��5�HH���  �'��u��5�HH���  ���uš�5�HH���  S�ҋȃ��E��t�W�t  ��5�HH���   h�  S3��҃����  ���_�u����    ��5�Hl�U�B�IWP�ы�������   ��5�F�J\�UP�A,R�Ѓ���t�K�Q�M�  ��5�F�J\�UP�A,R�Ѓ���t�K�Q�M�l  �E��;Pt&�F��5�Q\�J,P�EP�у���t	�MS�<  ��5�v�B\�M�P,VQ�҃���t�M�CP�  ��5�QH�E����   �E�h�  PG���у�;�����_^�   [��]� ��������U�조5�HH���   ]�������������̡�5�PH���   Q��Y��������������U�조5�HH���  ]��������������U�조5��P���   V�uW�}���$V�����E������At���E������z����؋�5�Q�B,���$V����_^]����������������U���0�5�U�V�u�U��]�W�P�}���   �E�PV�M�Q����� �@�@�E�����E��Au�����������z���������������z�����������Au������������z)���١�5�]��ɋ��]��]��P�RH�E�PV��_^��]���������Au������������������U�조5�HH�]��U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�HH�h�  �҃�������������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�HH�Vh  �ҋ�������   �EPh�  �0%  ����t]��5�QHj P���   V�ЋMQh(  �%  ����t3��5�JH���   j PV�ҡ�5���   �B��j j���Ћ�^]á�5�H@�QV�҃�3�^]�������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�HH�Vh�  �ҋ�����u^]á�5�HH�U�E��  RPV�у���u��5�B@�HV�у�3���^]�������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�HH�I]�����������������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�PH�EPQ���  �у�]� �U�조5�PH�EPQ���  �у�]� ̡�5�PH���  Q�Ѓ�������������U�조5�HH���  ]��������������U�조5�E�HH�U0�E,R�U(P�E$R�U P�ER�U���\$�E�$P��P  R�Ѓ�,]������������̡�5�PH���  Q�Ѓ�������������U�조5�PH�EP�EPQ���  �у�]� ������������̡�5�PH��  Q�Ѓ�������������U�조5�PH�EP�EP�EPQ���  �у�]� ��������̡�5�PH���  Q�Ѓ������������̡�5�PH���  Q�Ѓ�������������U�조5�PH�EPQ��  �у�]� �U�조5�PH�EPQ��  �у�]� ̋������������������������������̡�5�HH���  ��U�조5�HH���  ]��������������U�조5�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ���������U�조5�PH�E0P�E,P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ���  �у�0]�, ��������̡�5�PH��,  Q�Ѓ�������������U�조5�PH�EPQ��X  �у�]� ̡�5�PH��\  Q�Ѓ�������������U�조5�HH��0  ]��������������U�조5��W���HH���   j h�  W�҃��} u�   _��]� Vh�  �  ��������   ��5�HH���   j VW�҃��M��S�  ��5�P�E�R0Ph�  �M����E��5�P�B,���$h�  �M��Ћ�5�Q@�J(j �E�PV�у��M��\�  ^�   _��]� ^3�_��]� �����U��S�]�; VW��u7��5�U�HH���   RW�Ѓ���u��5�QH���   jW�Ѓ���t�   �����   ��5�QH���   W�Ѓ��} u(��5�E�QH�M���  P�ESQ�MPQW�҃��B�u��t;��5�U�HH�ER�USP���  VRW�Ћ�5���   �B(�����Ћ���uŃ; u��5�QH���   W�Ѓ���t3���   �W��u1��5�QH���   �Ћ�5�E�QH���   PW�у�_^[]� ��5�BH���   �у��} u0��5�M�BH�U���  Q�Mj R�UQRW�Ѓ�_^��[]� ��5�QH�h  �Ћ؃���u_^[]� ��5���   �u�Bx���Ћ�5���   P�B|���Ѕ�tU��5�E�QH�MP�Ej Q���  VPW�у���t��5���   �ȋBHS�Ћ�5���   �B(���Ћ���u�_^��[]� ��������������U��EV���u��5�HH���  �'��u��5�HH���  ���u��5�HH���  V�҃���u3�^]� P�EP���N���^]� ���������U���D��5�HH���   S�]VWh�  S�ҋ�5�HH���   3�Wh�  S�u܉}��҃��E�}�}��}�;��>
  ��5���   �B���Ћ�5=�  �  �QH���   Wh:  S�Ћ�5�QH�E����   h�  S�Ћ�5�QHW�����   h�  S�uԉ}��Ћ�5�QH�E苂  S�Ћ�5�QH�EЋ��  S�Ѓ�(�E��E����~~�M���M�I �MЅ�tMj�W�х�����t@�@�Ẽ|� �4�~����%�������;�u/���P���;E�~�E؋�����E���E�;Pu�E���E��E�G;}�|��}� ��   �u�j S���  ����  ���  ��ti���=  �}�;�u^��5�H���  �4�h���h�  V�҃��E���b  �M��E��I  ��t�}� t��tVP�E�P�PU ����}܋�5�Q���  �4�h���h�  V�Ѓ��E����  �M�3�;�t;�tVQP� U ���E�;�~-��5�Qh���h�  P���   �Ѓ��E�;���  ��5�E��QH��  j�PS�у�����  �u�;�tjS���u  ���{  ���  �E���}��5�BH���   Wh�  S�у�3��E�}�9}��]  �}���}����$    �MЅ��J  �U�j�R躃������6  �M̍@�|� ���]�~����%�������9E���  ��������E�3�3ɉE܉M�9C��   ��$    �����������ti�]������������M�ҋ9�<��}�҉T��y�]��|��]��z�|��y�]��|��]��z�|��I�}��]��L��M��}ȃ��T����M�A�M�;K�v����E؅��0  �+U�j��PR�M��w�  �M�v���E�3�+��U��E��ʋE�;E���   �}� �U����E�t4�U�M��@���P�Q�P�Q�P�Q�P�Q�@�A�M��Eȍ@�E��Ћ��P�Q�P�Q�P�Q�P�Q�@�A;]�}_�UȋE�9�uT�ȋL�����������w0�$���U���4���M���t���U���t��	�M���t��M���;]�|��E܃�F�M�;]������U�;U��  �U�R�yj���E�P�pj���M�Q�gj����_^3�[��]Ë�M�3�;G�Å���   �E�v�ЋW��R�ы��Q�P�Q�P�Q�P�Q�P�I�H�O��I�M�ы�P�Q�P�Q�P �Q�P$�Q�P(�I�H,��@�E�ЋU�Lv�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��t8�G�U�@�ʋU�Lv	�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�G��w��U��@�ʋU�F�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A��w��U�F�@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�7F��t=�G�U��@�ʋU�v�ʋ��P�Q�P�Q�P�Q�P�Q�@�A�wF���O�E�@���E��}�;E�������U�R�\h���E�P�Sh�����  ���   �B����=  ��  ��5�QH���   j h(  S�Ћ�5�QH�����   h(  S�ЋЃ�3��U؅�~"��ǅ�t�|� t�4N��tN�@;�|�u��u܋�5�Q���  �4v�h���hK  V�Ѓ��E�����   �M��t��tVQP�O ���u؋�5�Q���  �h���hP  V�Ѓ��E���tP��t��tVWP��N ���M����+�5�RH��PQ�E���   S�Ѓ���u�M�Q�g���U�R�	g����_^3�[��]á�5�HH���   j h�  S�҉E���5�HH���   j h(  S��3�3���3��E��}ĉ]�9]��:  �U��څ��  �E�    ����   �U�<��v��   ����U��:��\:�Y�\:�Y�\:׉Y�Z�Y�R�Q�U��\�EԉY�\�T�Y�Z�Y �Z�Y$�Z�Y(�R�]��Q,�U�@����0��;�|��}ă|� �t   �U��M�ύI�ʋU�v���A�B�A�B�A�B�A�B�I�J�E���ЋE�Tv�Ћ��A�B�A�B�A�B�A�B�I�J�U���<ډ}�C�]�;]�������M�3�3�;�~�U���$    �t���   @;�|��U�R�Ge�����E�P�;e����_^�   [��]�[�e�p�{�������������U��E� �M+]� ���������������U��V��V�Ե��5�Hl�AR�Ѓ��Et	V�h������^]� ���������̋�� 8����������8����������̅�t��j�����̡�5�P��  �ࡰ5�P��(  ��U�조5�P��   ��V�E�P�ҋuP���:�  �M��r�  ��^��]� ��������̡�5�P��$  ��U�조5�H��  ]��������������U�조5�H���  ]�������������̡�5�H��  ��U�조5�H���  ]��������������U�조5�H��x  ]��������������U�조5�H��|  ]��������������U���EV���8�t	V�f������^]� �������������̸   � ��������� ������������̸   � �������̸   � �������̸   � �������̸   � ��������� �������������3�� �����������3�� �����������3�� �����������3�� �����������3�� �����������3�� ����������̸   � �������̸   � �������̸   � ��������U���   V�����  �����   �ESP�M��ȭ  ��5�Q�J�E�P�ы�5�B�Pj j��M�h<�Q�҃��E�P�M�茭  j j��M�Q�U�R��d���P�T�  ��P�M�Q臱  ��P�U�R�z�  ���P���  ���M������  �M�蹭  ��d���训  �M�覭  ��5�H�A�U�R�Ѓ��M�芭  ��[t	V��  ����^��]� ���U��EVP���a�  �����^]� �����Q���  Y���������U��E�M�U�H4�M�P �U��M�@���@8p��@<@7�@@���@D�6�@HP7�@L���@P 7�@l 7�@X���@\7�@``7�@d���@T�7�@h���@pP��@t`��P0�H(�@,    ]��������������U���   h�   ��`���j P�G �M�U�Ej Q�MRPQ��`���R�����E �Uh�   ��`���Q�E��ERPj�%�����8��]��������������̋�`<����������̋�`@����������̋�`����������̋�`����������̋�`4����������̋�`(����������̋�`����������̋�`,����������̡�5�H\�������U�조5�H\�AV�u�R�Ѓ��    ^]�������������̡�5�P\�BQ�Ѓ���������������̡�5�P\�BQ�Ѓ����������������U�조5�P\�EPQ�J�у�]� ����U�조5�P\�EP�EPQ�J�у�]� U�조5�P\�EPQ�J�у�]� ���̡�5�P\�BQ�Ѓ����������������U�조5�P\�EPQ�J �у�]� ����U�조5�P\�EP�EPQ�J$�у�]� U�조5�P\�EP�EP�EPQ�J(�у�]� ������������U�조5�P\�EPQ�J0�у�]� ����U�조5�P\�EPQ�J@�у�]� ����U�조5�P\�EPQ�JD�у�]� ����U�조5�P\�EPQ�JH�у�]� ���̡�5�P\�B4Q�Ѓ����������������U�조5�P\�EP�EPQ�J8�у�]� U�조5�P\�EPQ�J<�у�]� ����U���SVW�}��j �ωu���  ��5�H\�QV�҃���S����  3���~=��I ��5�H\�U�R�U��EP�A(VR�ЋM��Q���X�  �U�R���M�  F;�|�_^[��]� ���������������U���VW�}�E��P��蘿  �}� ��   ��5�Q\�BV�Ѓ��M�Q���q�  �E���t]S3ۅ�~H�I �UR���U�  �E�P���J�  �E;E�!����5�Q\P�BV�ЋE@���E;E�~�C;]�|�[_�   ^��]� _�   ^��]� � �������������U���d�}W��t�   _��]� ���Pt�U�S�U�]�]�S�҉E��u[�   _��]� ��5�U�HH��   VRS�Ћ�5�Qd�J<�E��EP�эU�j/R�������E�jP�ק����5�Qd�E�JpVSP�у�(3�j ��u��5�Bd�U�@�M�QR�����5�Qd�M�R�E�PQ��3���9u~a3�;u���;�uO�E��RxVP�M�Q����� �U��@�]��@�]��������t��5�Hd�E���   j j�U�RP�у�F;u|�C���W���^[�   _��]� �������U����E�P�P�]� �������������  �������������3�� �����������U����   �ES��t
���[��]� ��5�PH�M�R,VW��$���P�ҋ���Pt�   �}��}W���E�����3��҅���   ���PxVW�M�Q����� �@�@���������A�|   �E���5�ˋUR�U��E����M����E������]��E����E��E������E������]��E������E��E������E������]�Hd�E�IP�ERP�у���t�E�u�t������؋�BtW��F��;��A����E�_^[��]� �����U�����5SVW�}��H@�Q8j W�ҋ]��Rx��SW�M�Q���ҋE�@��E�R|�Ƀ��ɋ�� �@0�E��������@H�E��������@ ���@�@8�����@P�����@(�����@�@@�����@X����S����������X�X�EP��_^�   [��]� ���������3�� �����������3�� ����������̸   �$ ��������� �������������� �������������� �������������3�� �����������3�� �����������U��UP�EQWRPV���������   ǆ�   �ǆ�   p7ǆ�   �6ǆ�   ��ǆ�   0�ǆ�   07ǆ�   ��]������������U�조5�P�B<��   V�u���Ѕ�t�Mj VQ���������u^��]�SWh   ������j R��= �]�E�}�M SP3��������(������E�@���t�E� ��� t�E� ���y�E�О_��[t�E���U�Eh   ������QRPj貟����^��]����������̋�`\����������̋�`l����������̋�`P����������̋�``����������̋�`p����������̋�`D����������̋�`d����������̋�`X����������̋�`h����������̡�5�PD�BQ�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�BQ�Ѓ����������������U�조5�PX��Q�
�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ���������U�조5�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�조5�PX��Q�J�E�P�ыM���P�Q�P�Q�P�Q�P�@�Q�A������]� ��������U�조5�PX��`VWQ�J�E�P�ы��E���   ���_^��]� �������������U�조5�PX�EPQ�J�у�]� ����U�조5�PX�EPQ�J�у�]� ����U�조5�PX�EPQ�J�у�]� ����U�조5�PX�EPQ�J�у�]� ����U�조5�PX�EPQ�J$�у�]� ����U�조5�PX�EPQ�J �у�]� ����U�조5�PD�EP�EPQ�J�у�]� U�조5�HD�U�j R�Ѓ�]�������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�HD�	]��U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�HD�U�j R�Ѓ�]�������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�U�HD�Rh2  �Ѓ�]����U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�U�HD�RhO  �Ѓ�]����U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�U�HD�Rh'  �Ѓ�]����U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�HD�j h�  �҃�����������U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�HD�j h:  �҃�����������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U���3��E��E���5���   �R�E�Pj�����#E���]�̡�5�HD�j h�F �҃�����������U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�HD�j h�_ �҃�����������U�조5�H@�AV�u�R�Ѓ��    ^]��������������U��E����u��]� �E���5�E�    ���   �R�E�Pj������؋�]� ̡�5�PD�B$Q�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ���������������̡�5�PD�B(Q�Ѓ���������������̡�5�PD�BQ�Ѓ����������������U���V�u�W�}�������Dz�F�G������D{:�G����$�f: �F��$�]��V: �E���������D{_�   ^��]�_3�^��]���������������������U���VW�M��`�  �E�}��t-��5�Q4P�B�Ѓ��M��u蘏  _3�^��]Ë�R(���5�H0�QW�҃��M��tԋ�R Q�MQ���ҋ�5�P�B �M��Ѓ��t��5�Q0�Jx�E�PW�у��M��.�  _��^��]�������U�조5�P�B VW�}�����=NIVb��   ��   =TCAbtR=$'  t6=MicM��   ��5�Q���   j hIicM���ЋWP�B����_^]� ��BW����_�   ^]� ��5�Q���   j hdiem���ЋWP�B����_^]� =INIb��   �~ u���B���F   ��_^]� �~ t���B����_^]� =atniDt5=ckhct=ytsdu?��B����_�F    3�^]� ��B����_^]� �A���_3�^]� =cnys����_3�^]� ������V���L���5�H0�Vh ��҉F���F    ��^�����V��F�L���t��5�Q0P�B�Ѓ��F    ^�����̡�5�P0�A���   P�у����������U�조5�P0�E�I���   PQ�҃�]� �������������̡�5�I�P0���   Q�Ѓ���������̡�5�P0�A���   j j j j j j j j j4P�у�(������̡�5�P0�A���   j j j j j j j j j;P�у�(�������U�조5�P0�E�IPQ���   �у�]� ��������������U����E V��P�M��;�  ��5�E�Q�R4Ph8kds�M��ҡ�5�E     �H0���   �U R�U�E�P�Ej R�UP�ER�UP�FRj2P�ыu ��(�M����  ��^��]� ��������������̡�5�I�P0���   Q�Ѓ����������U��V��F��u^]� ��5�Q0�M ���   j j j j j Q�Mj QjP�ҡ�5�H0�U�E���   R�UP�ER�UP�Fj RP�у�D^]� ���̋A��uË�5�Q0P�B�Ѓ������̋A��u� ��5�Q0P�B�Ѓ�� �U��Q����u�E�    �P��]� �E�H� V�5�5�v0Q�MQP���   R�U�R�Ћu�    �F    ��5���   j P�BV�Ћ�5���   �
�E�P�у�$��^��]� �������U�조5�P0�E�I�RPQ�҃�]� �U��A��t)��5�Q0�M���   j j j j j j Qj jP�҃�(]� ���������U��Q��u3�]� �E�H� V�5�5�v0Q�MQPR�V�҃�^]� ����������U��Q��u3�]� �E�H� V�5�5�v0QP���   R�Ѓ�^]� �����������U��Q��u3�]� �E�H� V�5�5�v0Q�MQPR�V\�҃�^]� ����������U��y u3�]� V�u�W�}�؉��ډ��5�P4�A�JhWVP�ы�ډ����ى_^]� �����U��A��u]� ��5�Q4�M�RhQ�MQP�҃�]� ����U��A��u]� ��5�Q4�M�RpQ�MQP�҃�]� ����U��y u3�]� V�u�W�}�؉��ډ��5�P4�A�JpWVP�ы�ډ����ى_^]� �����U���$VW��htniv�M��	�  ��5�P�E�R4Phulav�M��ҡ�5�P�B4hgnlfhtmrf�M��Ћ�5�E�Q�R4Phinim�M��ҡ�5�P�E�R4Phixam�M��ҡ�5�P�E�R4Phpets�M��ҡ�5�P�E�R4Phsirt�M��ҋE �}$=  �u�����t.��5�QP�B4h2nim�M��Ћ�5�Q�B4Wh2xam�M��ЋU�M�QR�E�P���K�����5���   P�B8�Ћ�5���   �
���E�P�у��M��(�  _��^��]�  ��������������U���$V��htlfv�M�躆  �E��5�P�B,���$hulav�M��Ћ�5�E,�Q�R4Phtmrf�M����E��5�P�B,���$hinim�M����E��5�Q�B,���$hixam�M����E$��5�Q�B,���$hpets�M��Ћ�5�ED�Q�R4Phsirt�M����E0��������������Dzw�E8������Dzm�؋�5�E@�Q�R4Phdauq�M��ҋM�E�PQ�U�R���������5���   P�B8�Ћ�5���   �
���E�P�у��M��ʅ  ��^��]�@ �ء�5�P�B,���$h2nim�M����E8��5�Q�B,���$h2xam�M����V���U���$V��hgnrs�M��*�  �E��5�E��E�   �Q���   �E�Pj�M��ҡ�5���   ��U�R�ЋM��5�M����E�   �B���   �M�Qj�M��ҡ�5���   ��U�R�ЋU���M�QR�E�P���������5���   P�B8�Ћ�5���   �
���E�P�у��M�誄  ��^��]� �U���$V��hCITb�M��J�  ��5�P�E�R8PhCITb�M��ҡ�5�P�E�R4Phsirt�M��ҡ�5�P�E�R4Phulav�M��ҋM�E�PQ�U�R��������5���   P�B8�Ћ�5���   �
���E�P�у��M����  ��^��]� U��E��Vj ��P�M�Q�M��  �UPR���)�����5�H�A�U�R�Ѓ���^��]� ����������U��E,��UPj ���T$�$htemf�E$�� �\$�E�\$�E�\$�E�$R�O���]�( �����������U��E,��Pj ���T$�U�$hrgdf�E$�� �б���@������\$�E�����\$�M���\$�E�$R�����]�( ���U��E,��Pj ���T$�U�$htcpf�E$�� �p������\$�E���\$�}�\$�E�$R����]�( ���������������U��Q��u3�]� �E�E�H� V�5�5�v0Q�M Q�M���\$�E�$QPR�V(�҃�$^]� ������U��Q��u3�]� �E�H� V�5�5�v0Q�MQPR�V,�ҋU3Ƀ�9M^���
]� �������������U��Q��u3�]� �E�H� V�5�5�v0Q�MQPR�V,�҃�^]� ����������U��Q��u3�]� �E�H� V�5�5�v0Q�MQPR�V0�҃�^]� ����������U��SVW���W��t$�E�H�5�5�^0� �uQVP�C0R�Ѓ���u	_^3�[]� �W��t��E�H� ��5�[0Q�NQPR�S0�҃���t̋W��tŋE�H� �=�5�0Q��VP�G0R�Ѓ���t�_^�   []� ��U��Q��u3�]� �E�H� V�5�5�v0Q�MQ�MQPR�V<�҃�^]� ������U��QV3�W��u3��,�E�H� �5�5�v0Q�MQPR�V,��3Ƀ�9M�������5�M�B�P0VQ�M�ҋ�_^]� ����U��AV��u3��"�M�Q�	�5�5�v0R�URQP�F,�Ѓ�����5�Q�E�M�R4PQ�M�ҋ�^]� ���������������U��A��V��u3��"�M�Q�	�5�5�v0R�U�RQP�F0�Ѓ�����5�E��Q�E�M�R,���$P�ҋ�^��]� �����U�����V���U��V�U��]�W��t$�E�H� �=�5�0Q�M�QPR�W0�҃���u
_3�^��]� �V��t�E�H� �=�5�0Q�M�QPR�W0�҃���tˋV��tċE�H� �5�5�v0Q�M�QPR�V0�҃���t���5�P�M�RH�E�PQ�M��_�   ^��]� �����������U��� ��A�U�V�U�W�]���u3��&�M�Q�	�5�5�v0R�U�R�U�RQP�F<�Ѓ����E�}���t��5�Q�RH�M�QP���ҋE���t��5�E��Q���$P�B,����_��^��]� U�조5�P�E���   Vj ��MP�ҋM$�U Q�MR�Uj Q�MR�UQPR���o���^]�  ����������U�조5��P�E���   V���$��MP���E8�E@�M,�Uj P���\$�E0�$Q�E$�� �\$���E�\$�E�\$�$R�K���^]�< ������U�조5��P�E���   V���$��MP����Ej j ���T$���$htemf�E$�� �\$�E�\$�E�\$�$P�����^]�$ �����������U�조5��P�E���   V���$��MP����j j ���T$�E�$hrgdf�E$�� �б�����@������\$�E�����\$�M���\$�$P�X���^]�$ ���U�조5��P�E���   V���$��MP����j j ���T$�E�$htcpf�E$�� �p��������\$�E���\$�}�\$�$P�����^]�$ ���������������U�조5��0V��H�A�U�WR�Ћ�5�Q�M���   ���E�PQ�M�E�P�ҋ���5�H�A�U�R�Ћ�5�Q�J�E�PW�ы�5�B�P�M�Q�ҋE�U��Pj �M�QR��������5�H�A�U�R�Ћ�5�Q�J�E�P�у�_��^��]� U���dV��M�蟃  ��5�Q���   P�EP�M�Q�M��P�M��)�  �M��a�  j j �E�P�M���  �MPQ���%�����5���B�P�M�Q�҃��M��&�  �M���  ��^��]� �����U���P��EV�]���W�}����t��5�Q���$P���   �����]����5�U��UЍE��]ȋQ�M���   PQ�E�P���ҋ�M��P�U�H�M�P�U�H�M��P�F�U��u_^��]� �M�E�Q�	�5�5�v0R�U R���\$�U��E��$RQP�F(�Ѓ�$_^��]� ���������������U���0�E�M���u��5�H���   �҅�u��]� SVW���Z  ��htlfv�MЉu�*y  �E�}��5�X�U�����$�# �]��G�$�# �}�S,�M��$hulav�ҡ�5�P�B4hmrffhtmrf�M��Ћ}���5�M�Y���$�E# �]��G�$�7# �}�S,�M��$hinim�ҋ}���5�M�X���$�	# �]��G�$��" �}�S,�M��$hixam���衰5�P�B,���$hpets�M��Ћ�5�Q�B4j hdauq�M��Ћ�5�Q�B4Vhspff�M��Ћ�5�E �Q�R4Phsirt�M��ҋM�E�PQ�M��U�R������5���   P�B8�Ћ�5���   �
���E�P�у��M���w  _��^[��]� U��E��V���u��5�H���   �҅�u^��]� ���X  �E�F��u3��"�M�Q�	�5�5�v0R�U�RQP�F0�Ѓ����E���x��M������\$�M��$�l�  ��M��P�Q�P�Q�@�A��^��]� ����������U���0�5�]�V���M�]�P���   �E�PQ�M�E�P�ҋ�P�M��Hj �U�P�E P�M��MQ�M�U��UR�U�E�PQR������^��]� ���������������U�����UV�]���E�P�]��ERP������5�Q�M�R@���E�PQ�M�ҋ�^��]� ����������U��A��u]� �M�Q�	V�5�5�v0Rj j j j j j Qj1P���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��A��u]� ��5�Q0�M���   j j j j j j j Qj-P�҃�(]� �����U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j j Q�MQj j j)P�ҋE���(��]� ��U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�Mj Qj j j)P�ҋE���(��]� ��U��A��u]� ��5�Q0�M���   j j j Q�MQ�MQ�Mj Qj/P�҃�(]� ���������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj'P�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQj,P�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�MQ�MQjP�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�MQ�MQjP�ҋE���(��]� ����������U�조5�P0�E�I���   j j j P�EP�EP�Ej Pj.Q�҃�(]� ��������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj:P�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj*P�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj	P�ҋE���(��]� ��������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj Qj
P�ҋE���(��]� ��������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��A��u]� ��5�Q0�M���   j j j Q�MQ�MQ�Mj QjP�҃�(]� ���������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj QjP�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj Q�MQ�MQ�MQ�Mj Qj>P�ҋE���(��]� ������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� �M�Q�	V�5�5�v0R�Uj j j j R�URQjP���   �Ѓ�(^]� �����������U����ESVW�M�P�M���  �MQ�U�R�M��X�  ��tm�}��E��tN��5���   P�BH�ЋM��I����tQ�W�7��5�[0R�U�j j j j RP���   VjQ�Ѓ�(��t"�MQ�U�R�M���  ��u�_^�   [��]� _^3�[��]� ��������������U��A��u]� �M�Q�	V�5�5�v0Rj j j j j j QjP���   �Ѓ�(^]� ���������������U��Q�A��u��]� ��5�E�    �Q0���   �M�Q�Mj j Q�MQ�MQ�Mj QjP�ҋE���(��]� ��������������U��A��u]� ��5�Q0�M�RDQ�MQ�MQP�҃�]� U��A��u]� ��5�Q0�M�RHQ�MQ�MQ�MQ�MQ�MQP�҃�]� ���̋A��uË�5�Q0P�BX�Ѓ�������U��A��u]� ��5�Q0�M�RLQ�MQP�҃�]� ����U��A��u]� ��5�Q0�M�RP��   �QP�҃�]� ��U��A��u]� ��5�Q0�M�RPQP�҃�]� ��������U��A��u]� ��5�Q0�M�RTQ�MQ�MQ�MQP�҃�]� ������������U�조5V�u�VW���H4�R�ЋE�F    �~�H� ��5�R0Q�MQ���   VP�GP�у�3҅��F_^��]� ���U��A��u]� ��5�Q0�M���   j j j j j Qj j jP�҃�(]� �����U��E��u]� �@    �@�I��5�R0P�EPQ���   �у�]� ������̡�5�I�P0���   j j j j j j j j j0Q�Ѓ�(�������U��E��u��5� ��5�R0�I�R@V�uVP�EPQ�҃�^]� �����������U�조5�P0�E�I�RdP�EP�EP�EP�EPQ�҃�]� �U�조5�P0�E�I�RpP�EP�EP�EP�EPQ�҃�]� �U��E�P� V�5�5�v0R�UR�UR�UR�URP�A�NhP�у�^]� ��������U��E� ��5�R0j j j j j j j P�A���   jP�у�(]� �����������U��E� ��5�R0j j j j j jj P�A���   jP�у�(]� �����������U��E� ��5�R0j j j j j j j P�A���   jP�у�(]� �����������U���V��M��Og  �E�H� ��5�R0Q�M�Q���   j j j j j P�Fj8P�ы���(��t�M�U�R�{g  �M��cg  ��^��]� ����������U��E�P� V�5�5�v0R�URj j j j j P�A���   j9P�у�(^]� �����U��E�P� V�5�5�v0Rj j j j j j P�A���   j"P�у�(^]� �������U��E�P� V�5�5�v0Rj j j j j j P�A���   j5P�у�(^]� �������U��E�P� V�5�5�v0R�Uj j j j Rj P�A���   j<P�у�(^]� �����U�조5�P0�E�I���   j j P�EP�EP�EP�Ej Pj3Q�҃�(]� ������U�조5�UVj j j j j R��H0�E�Vj P���   jR�Ћ�5�Q0�E�N�RtPQ�҃�0^]� ��U�조5�P0�E�I���   j j j j j j Pj jQ�҃�(]� �������������̡�5�P0�A���   j j j j j j j j jP�у�(�������U�조5�P0�E�I���   j j j j j j j PjQ�҃�(]� �������������̡�5�P0�A���   j j j j j j j j j(P�у�(�������U�조5�P0�E�I���   j j j j j j P�EPj&Q�҃�(]� ������������U�조5�P0�E�I���   j j j j P�EP�Ej Pj+Q�҃�(]� ���������̡�5�P0�A���   j j j j j j j j jP�у�(������̡�5�P0�A���   j j j j j j j j j#P�у�(�������U��QS�]VW�}�M���t��5�P���   j j���Љ�u��t��5�Q���   j j���Љ��5�Q0�E��H�R`VWQ�҃�_^[��]� �U�조5�P0�E�I���   P�EP�EPQ�҃�]� �����̡�5�P0�A���   j j j j j j j j j P�у�(������̸   ����������̸   ��������������������������̸   � ��������3�� �����������3���������������� �������������V���L���5�H0�Vh ��҉F3��F�F������F   ��^�������V��F�L���t��5�Q0P�B�Ѓ��F    ^������U��V��F�F    ��tn��5�Q0j j j j j j j j jP���   �Ћ�5�Q0�E�MP�E���   Q�MP3�9EQ�N��j ��
PQ�҃�D��t�~ t
�   ^]� 3�^]� �������U��E�A�I��u3�]� ��5�B0Q�H�у�]� ����U�조5�P�B S�]V�����=ckhc��   ��   =cksate=TCAb��   ��5�Q���   Wj hdiem���Ћ���BSW���F   �Ѓ~ ��t��t��u3Ƀ���Q���C���_^��[]� �~ tn��B����^[]� �~ tY��5�Q0�F���   j j j j j j j j j P�у�(��t+�F    ^�   []� =atnit�URS���l���^[]� ^3�[]� ��������������U��V��~ ��   W�}����   �$�x��E;E��   �r�M;M��   �d�U;U��   �V�E;E��   �H�E;E~@;E��   �5�E;E|-;E~v�&�E;E|;E|g��E;E~;E~X��M;MuN��5�M�B0�V���   j j j j j j j QjR���E��(j���\$�E�$W��i�����F    _^]� ��������������������U��V��~ �  �E W�}�E����   �$������]������   �   ���]����A��   �   ���]����A��   �t���]������   �b�E������A��uP��������   �E�E��������u3������A{}�,�E���������E������A�����E������DzU����ء�5�U�H0�F���   j j j j j j j RjP���E �U(��(R���\$�E�$W�h�����F    _^]�$ ���������5�N�Z�f�������������U���E �E�Uj���\$�E�\$�E�$PR�w���]�  ���U���E �E�Uj���\$�E�\$�E�$PR�G���]�  ���U���E �E�Uj���\$�E�\$�E�$PR����]�  ��̋�3�� ���H�H�H�������������VW��3����9~u��5�H4�V�R�Ѓ��~�~_^����U�조5�P4�E�I�RtPQ�҃�]� �U��U��t3�A��5�I0R���   P�ҋ�5�Q0�M���   QP�҃�]� ��5�P0�E�I�R|PQ�҃�]� ������̡�5�P4�A�JP�у������������̡�5�P4�A�JP�у������������̡�5�P4�A�JP�у������������̡�5�P4�A�J|P�у������������̡�5�P4�A���   P�у����������U�조5�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�조5�P4�E�I�RP�EP�EP�EPQ�҃�]� �����U�조5�P4�E�I�R PQ�҃�]� �U�조5�P4�E�I�R$PQ�҃�]� �U�조5�P0�E�I���   P�EP�EP�EPQ�҃�]� ��U�조5�P4�E�I���   PQ�҃�]� ��������������U�조5�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�조5�P4�E�I���   P�EP�EP�EP�EPQ�҃�]� ��������������U�조5�P4�E�I�R(PQ�҃�]� �U�조5�P4�E�I�R,P�EP�EPQ�҃�]� ���������U�조5�P4�E�I�R0P�EPQ�҃�]� ������������̡�5�P4�A�J4P��Y��������������U���S�]V3����5W�~�E�E��QP���   j���Ћ�5�E��Q���   j j���Ћ�5�E�Q0�EP�G�M�Q�J`P�ы�5�B4�N�PQ�ҋ�5�Q0�Rhj �M�Q�M�Q�M�Q�M�QP�F�HQ�҃�,�} _^[t(�} t(�E��M�;�~<�U��;�}3�E�M�;�~)�U���} u�E��M�;�~�U��;�}�   ��]� 3���]� U�조5�P4�E�I�R8PQ�҃�]� �U�조5�P4�E�I�R<PQ�҃�]� �U�조5�P4�E�I���   P�EPQ�҃�]� ���������̡�5�P4�A�J@P�у�������������U�조5�P4�E�I�RDP�EPQ�҃�]� �������������U�조5�P4�E�I�RHP�EPQ�҃�]� �������������U�조5�P4�E�I�RLP�EPQ�҃�]� �������������U�조5�P4�E�I�RPP�EPQ�҃�]� �������������U�조5SV�uW�����   �QV�҃�����   ��5���   �]�QS�҃�S��uA��5���   �Q@�ҋء�5���   �Q@V�ҋ�5�Q4�JPSP�GP�у�_^[]� ��5���   �H�у���uD��5���   �H8S�ы�5�؋��   �H@V�ы�5�J4�WSP�AHR�Ѓ�_^[]� hضh}  ��   ��5���   �BV�Ѓ�����   ��5���   �]�BS�Ѓ�S��uC��5���   �B@�Ћ�5���   �؋B8V�Ћ�5�Q4�JLSP�GP�у�_^[]� ��5���   �H�у���uD��5���   �H8S�ы�5�؋��   �H8V�ы�5�J4�WSP�ADR�Ѓ�_^[]� hضh�  �
hضh�  ��5�Q��0  �Ѓ�_^[]� �U�조5�P4�E�I��  P�EP�EP�EPQ�҃�]� ��U�조5�P4�E,P�E(P�E$P�E �IP�E�RTP�EP�EP�EP�EP�EPQ�҃�,]�( �������������U�조5�P4�E�I�RXP�EP�EP�EPQ�҃�]� ����̡�5�P4�A�J`P��Y�������������̡�5�P4�A�JdP�у�������������U�조5�P4�E�I��   P�EP�EP�EPQ�҃�]� ��U�조5�P4�E�I�R\P�EP�EP�EP�EP�EPQ�҃�]� �������������U�조5�P4�E�I�RhP�EPQ�҃�]� �������������U��V�uW��t��؉�}��t��ډ��5�P4�A�JhWVP�у���t��ډ��t��ى_^]� �U��V�uW��t��؉�}��t��ډ��5�P4�A�JpWVP�у���t��ډ��t��ى_^]� �U�조5�P4�E�I�RpP�EPQ�҃�]� �������������U���,V��~ ��   ��5�V�H4�AR�Ѓ} t ��5�Q0�RlP�F�HQ�҃�^��]� ��hARDb�MԉE��E�    �|R  P�M�Q�N�U�R������5���   ��U�R�Ѓ��M��R  ^��]� ������U�조5�P4�E�I�RlPQ�҃��   ]� ������������U�조5�E�P4�E�I���   P�E���\$�E�$PQ�҃�]� ����������U�조5�P4�E�I���   P�EP�EPQ�҃�]� �����̡�5�P4�A���   P�у���������̸   ����������̸   �����������U�조5V��H4�V�A$h�  R�Ћ�5�Q4�E�MP�EQ�MP�FQ�JP�у�2�^]� ��������U��U��@R�UR�UR�UR��]� �̸   � ��������3�� ������������ �������������3�� ������������ �������������U�조5�P4�E�I�RxP�EP�EP�EPQ�҃�]� �����U�조5�P0�E�I�I���   P�EP�EPQ�҃�]� ���U��QS�]VW�}�M���t��5�P���   j j���Љ�u��t��5�Q���   j j���Љ��5�Q4�E��H�RpVWQ�҃�_^[��]� �U��Q��5�P�B SVW�}���3���=INIb�/  �  =SACbvt+=$'  t
=MicM�  ��B$W����_�   ^��[��]� ��R3��E��E�EP�M�Q���҅�t��5�U�H4�E�R�VP�AR�Ѓ�_�   ^��[��]� =ARDb�  ��5�Q���   j j���Ћ�5�Qj �؋��   j���Ћ�5�Qj �E����   j���Ћ�5�Qj �E���   j���ЋM���RWP�EPQS����_�   ^��[��]� ��P����_�   ^��[��]� =NIVbetJ=NPIbt0=ISIbu\�>���)���P������P�G����_�   ^��[��]� ��BW����_^[��]� ��B����_�   ^��[��]� =cnyst_^��[��]� ��5�Q���   j hIicM���ЋWP�B ����_^[��]� �������������U�조5�P4�E�I�RTh����h����h����P�EP�Eh����h����h����h����PQ�҃�,]� ������U���V��hYALf�M��ZM  ��5�Q4�JlP�FP�у��M��|M  ^��]��������V���L���5�H0�Vh ��҉F���F    � ��F   ��^��������V��F�L���t��5�Q0P�B�Ѓ��F    ^������U�조5�P�B VW�}�����=cksat`=ckhct�MQW��譽��_^]� �Nj j j j j j �F   ��5�B0���   j j j Q�҃�(��t'_�F    �   ^]� �~ t��P����_^]� _3�^]� ���U�조5�H���  ]��������������U�조5�H0���   ]��������������U�조5�H0�U�E��VWRP���   �U�R�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�_��^��]������������U�조5�H0���   ]��������������U�조5�H0���   ]��������������U��Ej0P�P����]��������������U��Ej0P��k����P�P����]�����U��E�M��j0PQ�U�R��k����P�^P����5�H�A�U�R�Ѓ���]�������U��E�M�U��j0PQR�E�P��l����P�P����5�Q�J�E�P�у���]��U��Ej$P��O��3Ƀ�������]����U��Ej$P�k����P��O��3Ƀ�������]�����������U��E�M��Vj$PQ�U�R��j����P�O����53Ƀ��B�P����M�Q�҃���^��]��������U��E�M�U��Vj$PQR�E�P�l����P�9O����53Ƀ��B�P����M�Q�҃���^��]����U�조5�H�U�E���   RPj �у�]���������������U�조5�H�U�ER�UP���   Rj �Ѓ�]�����������U�조5�P4�E�I�R,P�EP�EPQ�҃�]� ���������U�조5�P4�E�I�R0P�EPQ�҃�]� ������������̡�5�P4�A�J4P��Y��������������U�����5�P���   VW�}j ��j���Ћ�5�E��Q���   j j���Ћ�5�E�Q0�EP�F�M�Q�J`P�ы�5�J0�E�P� R�U�R�U�R�U�R�U�R�VP�AhR�Ѓ�(�} _^t&�} t&�E��M�;�~8M�;�}1�E�M�;�~'M���} u�E��M�;�~M�;�}�   ��]� 3���]� ���������������U��ESVW�؅�u�Y��5�P�}���   j hdiuM���Ћ���tK;3u	_^3�[]� ��5�Q���   j hIicM����;�u��5�Q���   j h1icM���Шu��3_^�   []� �����U�조5�P�BT��(V�uhfnic���Ѕ�t��5�Q�ȋ��   j
�Ѕ���   ��5�Q�RPhfnic�E�P����P�M���F  �M���F  �u�E�P����F  �M���F  ��5�Q�B ���Ѓ��t��5�Q�B ���Ѕ�u��5�Q�B$hfnic���Ћ�5�E�Q�R8Pj
����^��]���������U�조5�P0�E�IP�EP�EP�EPQ���   �у�]� ��U�조5�P0�E�IV�p� ���   V�uj j j V�uVj Pj=Q�҃�(^]� ����U�조5�P0�E�IV�p� ���   V�uV�uj j j�Vj Pj=Q�҃�(^]� ���̡�5�I�P0���   j j j j j j j j j6Q�Ѓ�(�������U��V���L���5�H0�WVh ��ҋ}�F�E�F    �F   �L��F��5�Q���   ��j hmyal���ЉF��t��t�F    ��5�Q���   j
hhfed���ЉF_��^]� �����������U�조5�P�B VW�}�����=ytsdt�MQW�������_^]� ��5�B0�N���   Q�ҋ�P������_�   ^]� ��3���������������3�������������������������������3���������������3���������������3���������������3�� �����������U��V���PD�҅�t�E9Ft�F��PH����^]� �����̋A������������̋A��uË ��������������������̸�������������U���E�Y(]� ���U���(V���P(�M�Q���ҋN��t&��5�R0j j j j j j P���   j jQ�Ѓ�(��5�Q�J�E�P�ы�5�B�P�M�Q�ҋF����t ��5�Q0�RHj �M�Qj jj?j P�҃���5�H�A�U�WR�Ћ�5�Q�J�E�P�ыF����u3��;��5�E�    �J0�U�Rj j j h  
 j�U�Rh�  jP���   �Ћ}���(��5�Q�J�E�P�у���_u3�^��]Ë�5�B�P�M�Q�ҋF����t ��5�Q0�RHj �M�Qj j j8j P�҃���5�H�A�U�R�ЋF����t��5�Q0jP�BP�Ѓ���5�Q�J�E�P�у��M��A  Ph   h  K j;�U�Rh	��h�  ���w�����5�H�A�U�R�Ѓ��M���A  �F��t��5�Q0P�BX�Ѓ��F��t��5�Q0P�BX�Ѓ��F��t'��5�Q0j j j j j jj j jP���   �Ѓ�(j�v$�QF�����   ^��]�����U���SVW��j�N�K�  ��V�^(3ۉ^4�^8�^<��5�H0�Ah�   R�Ћ�5�Q�J�E�P�ы�5�B�PSj��M�h��Q�҃�SS�E�P�M�Q���E��  �]��+�����5�B�P�M�Q�҃�Sj�N苗  _^[��]����̍A�������������U��VW��~4 tA�I ��5�H��0  hضhj  ��j
�/O����5�HP�V �AR�Ѓ���uP9F4u�5�QP�Bh�N0�Ѓ~4 t<��5�Q��0  hضh�  �Ћ�5�QP�Bl���N0���n���_3�^]� �M�U�N8�V4��5�PP�Bl�N0�Ѓ~4 t%j
�N����5�QP�F �JP�у���u�9F4uۋ�5�BP�PhS�N0�ҋ^<�F<    ��5�PP�Bl�N0�Ћ�[_^]� ���U�조5�P�B ��@VW�}�����=MicMtI=fnic��   j�M���>  �uP���=?  �M��%?  ��5�Q�B4jj����_�   ^��]� ��5�Q���   j hIicM����=�����   htats�M��>  ��5�Q�B0j j�M��ЍM�Q�U�R�E�P���E��  �E�    茳����5���   �
�E�P�у��M��}>  �F�F   ��t��5�J0�QP�҃��EPW�������_^��]� ���������U��E��V��t3�^]� j�N�1�  j�
C���F    �v����t��5�H0�QV�҃��   ^]� ��������������j����  j�B����3�����������U��E3�h�����h  ���P�Ej BR�Uj PR�5���]� �U��Q�Q��u3���]� �E�H� V�5�5Q�M�Q�E�    �v0PR�V8�ҋ�����t@�E���t9��5�Q�M�RQP�ҋE�����t��5�QW��P�B��W������_��^��]� ������U�조5��V��H�A�U�R�ЋU���M�QR���D�������u��5�H�A�U�R�Ѓ�3�^��]� �M�Q�M�EG  ��5�B�P�M�Q�҃���^��]� �������U�조5��V��H�A�U�R�ЋU���M�QR��������M��5�P�R8�E�PQ�M�ҡ�5�H�A�U�R�Ѓ���^��]� �������������U���V��M��D  �M�E�PQ���������5���B�U�@<�M�Q�MR�ЍM��ME  ��^��]� ����U�조5�P�E���   Vj ��MP��h���h  �j j jj P�EP���#���^]� ��������������U�조5V�uW�����   �QV�҃�V��u,��5���   �Q@�ҋ�5�Q4�J P�GP�у�_^]� ��5���   �H�у���u.��5���   �H8V�ы�5�J4�WP�A$R�Ѓ�_^]� ��5�Q��0  hضh	  �Ѓ�_^]� �����U���4��5�H�QSVW�}W�ҡ�5�P�u���   ��3�SS�Ή]�Ћ�5�QS�E����   j���Ћ�;��L  �d$ �} ~l��5�Q�J�E�P�ы�5�B�Pj j��M�h��Q�ҡ�5�P�B<�����Ћ�5�Q�RLj�j��M�QP���ҡ�5�H�A�U�R�Ѓ���5�Q0�E����   VP�M�Q�ҋ�5�H�A�U�R�Ћ�5�Q�J�E�PV�ы�5�B�P�M�Q�ҡ�5�P�B<�����Ћ�5�Q�RLj�j��M�QP���ҡ�5�H�A�U�R�Ћ�5�Q�u���   �E��j ��
S���Ћ�5�Q���   �E�j �CP���ҋ����������_^[��]����������������U��E�PV��3Ƀ8������t�   3�h�����h  ���Pj AQj R�UR���M���^]� ��������U��E3҃8�@V�u ��V�uVR�UR�UR�UR�UPR����^]� ����������U��E�E43҃8��R�U<R�U(���\$�E,�$R�E �� �\$�E�\$�E�\$�@�E�$P����]�8 ��������������U��E�@3҃8��E��Rj ���T$�$htemf�E �� �\$�E�\$�E�\$�$P觰��]�  ���U��E�@3҃8��E��Rj ���T$�$hrgdf�E �� �б���@������\$�E�����\$�M���\$�$P�?���]�  �����������U��E�@3҃8��E��Rj ���T$�$htcpf�E �� �p������\$�E���\$�}�\$�$P�ۯ��]�  �������U��E3҃8��R�UR�UR�UR�UP�EPR����]� U��E3҃8V�u��V��RP�EP����^]� ����������U��Q��u3�]� �E�E�H� V�5�5�v0Q�M Q�M���\$���E�$QPR�V(�҃�$^]� ���U�조5�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U�조5�P�E���   Vj ��MP�ҋ���u�    �F^]� ��u9Ft�   ^]� ��������U�조5��P�E���   V���$��MP�ҋ���u�^�    ^]� ��u�F������D{�   ^]� ��^]� ����U���0�5�U�V�U���M�]�P���   �E�PQ�M�E�P�ҋ���̉�P�Q�P�Q�P�Q�P�@�Q�A���O	  ^��]� ��������U���0�5�]�S��V�]�W��P�M���   �E�PQ�M�E�P�ҋ�x�X��@�U��}�]��E����u�V�~�^_�    �F^[��]� ��u�E�P�NQ��������t�   _^[��]� ������������U���VW�}�M�;}us��5�P�u���   j htsem���Ѕ�uS��5�QP���   hrdem���Ѕ�u6�MQ�M�U�R�E�}�E��w�����t�E�M�P�  _�   ^��]� _3�^��]� U��SVW�}��;}u~��5�P�u���   j htsem���Ѕ�u^��5�QP���   hrdem���Ѕ�uA�M�E�A��t4��5�J0j �URWP�A,�Ѓ���t�MQ���  _^�   []� _^3�[]� ���������U���SVW�}��;}��   ��5�P�u���   j htsem���Ѕ�ug��5�QP���   hrdem���Ѕ�uJ�M��A�]���t;��5�J0j �U�RWP�A0�Ѓ���t�E������$�  _^�   [��]� _^3�[��]� �������U���4�ESW�}�M�;�t;Et	;E��   ��5�P�]���   j htsem���Ѕ���   ��5�QP���   hrdem���Ѕ�uj�M��U�U܉E��UԉE��]̉E�M�E�P�M�Q�M�U�U�R�E�P�}��1�����t+�E̋M�������E��X�E��X��  �   _[��]� _3�[��]� ��������U���SVW�}��;}��   ��5�P�u���   j htsem���Ѕ�uj��5�QP���   hrdem���Ѕ�uM��U�M��]���Q�M�]��E�R�E�P�}�������t%�E��������E��X�  �   _^[��]� _^3�[��]� ���̋A���X(Q�ȋB$��j j h����P8�����������������U�조5��@VW���H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�U���M�QR���   �M�Q�M�ҋ�5�H�A�U�R�Ћ�5�Q�J�E�PV�ы�5�B�P�M�Q�ҡ�5�H�I�U�R�E�P�ы�5�B�P�M�Q�ҡ�5�H�A�U�R�Ћ�5�Q�B����V�Ћ�5�Q�JV�E�P�у����  ��5�B�P�M�Q�҃�_^��]� ��U���SVW�}��;}��   ��5�P�u���   j htsem���Ѕ�ue��5�QP���   hrdem���Ѕ�uH��5�Q�J�E�P�ыM���U�R�E�P�}��E�    �]�����u ��5�Q�J�E�P�у�3�_^[��]� ��5�B�H����V�ы�5�B�P�M�VQ�҃����  ��5�H�A�U�R�Ѓ�_^�   [��]� ������U���V�u3ɍF��H�������5�M��M����   �RQ�M�QP�ҡ�5���   ��U�R�Ѓ���^��]� ����������U���\��5SV��H�A�U�WR�Ћ�5�Q�J3�Sj��E�h��P���F(�p��E��  �]��`�  ��5�JP�A(�U�R�Ћ�5�Q�J���E�P�ы�5�B�P�M�QW�ҡ�5�H�A�U�R�Ћ�5�Q�J�E�P�ы�5�B�@�M�Q�U�R�Ћ�5�Q�B<��8�M��Ћ�5�Q�RLj�j��M�QP�M���SS�E�P�M�Q���n�����5�B�P�M�Q�ҡ�5�H�A�U�R�Ћ�5�Q�J�E�P�у�htats�M��,  ��5�B�P0jj�M����F(��5�P�B,���$j�M��ЍM�Q�U�R�E�P���E��  �]��l�����5���   �
�E�P�у�9^4t[��5�BP�Ph�N0�ҋF4;�t�N8Q�Ѓ��F<�^8�^4���5�B��0  hضh�  �у���5�BP�Pl�N0�ҍM���+  _^[��]� ����U�����u�E�    �A]� ��u�Q;Ut�   ]� U�����u�E�    �Y]� ��u�A�E������D{�   ]� ���������U�����u�E�    �Y�E�Y�E�Y]� ��u3�A�E������Dz�A�E������Dz�A�E������D{�   ]� ���������������U��V�����u#�E�M�U�F�E�N�V�    �F^]� ��u�MQ�VR��������t�   ^]� �������������U��V��~ ���u��5�H4�V�R�Ѓ��E�F    �F    t	V���������^]� �������U��V��F�L���t��5�Q0P�B�Ѓ��E�F    t	V��������^]� ��������������U��V�����u �    ��5�H�A���UVR�Ѓ��#��u��5�Q�Rx�EP�N�҅�t�   ��5�H�A�UR�Ѓ�^]� ������̡�5�HL���   ��U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�HL�������U�조5�H@�AV�u�R�Ѓ��    ^]�������������̡�5�PL���   Q�Ѓ�������������U�조5�PL�EP�EPQ���   �у�]� �������������U�조5V��HL���   V�҃���u��5�U�HL���   j RV�Ѓ�^]� ��5���   �ȋBP�Ћ�5���   �MP�BH��^]� �����̡�5�PL��(  Q�Ѓ�������������U�조5�PL�EP�EPQ��,  �у�]� ������������̡�5�HL�Q�����U�조5�H@�AV�u�R�Ѓ��    ^]��������������U�조5�PL�E�R��VPQ�M�Q�ҋu��P���'  �M��'  ��^��]� ����U�조5�PL�EPQ���   �у�]� �U�조5�PL�EP�EPQ�J�у�]� ��5�PL�BQ�Ѓ���������������̡�5�PL�BQ�Ѓ���������������̡�5�PL�BQ�Ѓ����������������U�조5�PL�EP�EP�EPQ�J �у�]� ������������U�조5�PL�EPQ��4  �у�]� �U�조5�PL�EP�EP�EPQ�J$�у�]� ������������U�조5�PL�EP�EP�EP�EPQ�J(�у�]� �������̡�5�PL�B,Q�Ѓ���������������̡�5�PL�B0Q�Ѓ����������������U�조5�PL�EP�EPQ��  �у�]� ������������̡�5�PL���   Q�Ѓ�������������U�조5�PL�E��  ��VPQ�M�Q�ҋu��P���b%  �M��z%  ��^��]� ̡�5�PL�B4Q�Ѓ���������������̡�5�PL�B8j Q�Ѓ��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL���   ]��������������U�조5�PL�EPQ�J<�у�]� ���̡�5�PL�BQ��Y�U�조5�PL�EP�EPQ�J@�у�]� U�조5�PL�Ej PQ�JD�у�]� ��U�조5�PL�Ej PQ�JH�у�]� ��U�조5�PL�EjPQ�JD�у�]� ��U�조5�PL�EjPQ�JH�у�]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��]  W�M�Q�U�R���Ԁ  ���M�����O  ��t��5���   ��U�R�Ѓ�_^3�[��]Ë�5���   �J8�E�P�ы�5�����   ��M�Q�҃�_��^[��]��������������U���$3�V�E��E�E��P�M��E�   �E�   �E��  ��\  j�M�Q�U�R���=�  �M��EO  ��5���   ��U�R�Ѓ�^��]�����������U���$��5�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}��Z\  j�E�P�M�Q���  �M���N  ��5���   ��M�Q�҃�_^��]� ��U���$��5�UVW3���}܉}䋈�   �I(R�E�P�у��U�R�M��E��  �}��}���[  j�E�P�M�Q���9  �M��AN  ��5���   ��M�Q�҃�_^��]� ��U���$SVW3��E��P�M��}܉}��E��  �}��}��t[  W�M�Q�U�R���~  ���M�����M  ��t+�u���Y)  ��5���   ��U�R�Ѓ�_��^[��]� ��5���   �JL�E�P�ыu��P����)  ��5���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}��Z  W�M�Q�U�R����}  ���M����M  ��t+�u���(  ��5���   ��U�R�Ѓ�_��^[��]� ��5���   �JL�E�P�ыu��P���)  ��5���   ��M�Q�҃�_��^[��]� ���U���$SVW3��E��P�M��}܉}��E��  �}��}���Y  W�M�Q�U�R���4}  ���M����WL  _^��[t��5���   ��U�R�������]Ë�5���   �J<�E�P���]���5���   ��M�Q���E�����]���������������U���$SVW3��E��P�M��}܉}��E��  �}��}��DY  W�M�Q�U�R���|  ���M����K  ��t��5���   ��U�R�Ѓ�_^3�[��]Ë�5���   �J8�E�P�ы�5�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��X  W�M�Q�U�R����{  ���M�����J  ��t-��u��5����   ���^�U�R�Ѓ�_��^[��]� ��5���   �JP�E�P�ы�u�H��P�@�N��5�V���   �
�F�E�P�у�_��^[��]� �����̡�5�PL���   Q��Y��������������U�조5�PL�E���   ��jPQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U�조5�PL�E���   ��j PQ�M�Q�ҋM���P�Q�P�@�Q�A������]� �����������U���$SVW3��E��P�M��}܉}��E��  �}��}��W  W�M�Q�U�R���Dz  ���M����gI  ��t-��u��5����   ���^�U�R�Ѓ�_��^[��]� ��5���   �JP�E�P�ы�u�H��P�@�N��5�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��4V  W�M�Q�U�R���ty  ���M����H  ��t-��u��5����   ���^�U�R�Ѓ�_��^[��]� ��5���   �JP�E�P�ы�u�H��P�@�N��5�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��dU  W�M�Q�U�R���x  ���M�����G  ��t-��u��5����   ���^�U�R�Ѓ�_��^[��]� ��5���   �JP�E�P�ы�u�H��P�@�N��5�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}��T  W�M�Q�U�R����w  ���M�����F  ��t��5���   ��U�R�Ѓ�_^3�[��]Ë�5���   �J8�E�P�ы�5�����   ��M�Q�҃�_��^[��]��������������U����E3�V�]�E��E��E��P�M�E�   �E��  ��S  j�M�Q�UR���>w  �M�FF  ��5���   ��U�R�Ѓ�^��]� ���������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��oS  j�U�R�E�P����v  �M���E  ��5���   �
�E�P�у�^��]� ��������U���$��5�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���R  j�E�P�M�Q���Iv  �M��QE  ��5���   ��M�Q�҃�_^��]� ��U���$��5�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��jR  j�E�P�M�Q����u  �M���D  ��5���   ��M�Q�҃�_^��]� ��U���$��5�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}���Q  j�E�P�M�Q���Iu  �M��QD  ��5���   ��M�Q�҃�_^��]� ��U���$��5�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��jQ  j�E�P�M�Q����t  �M���C  ��5���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E���P  j�U�R�E�P���^t  �M��fC  ��5���   �
�E�P�у�^��]� ��������U���$SVW3��E��P�M��}܉}��E��  �}��}��P  W�M�Q�U�R����s  ���M�����B  ��t-��u��5����   ���^�U�R�Ѓ�_��^[��]� ��5���   �JP�E�P�ы�u�H��P�@�N��5�V���   �
�F�E�P�у�_��^[��]� ������U���$SVW3��E��P�M��}܉}��E��  �}��}���O  W�M�Q�U�R���s  ���M����'B  ��t��5���   ��U�R�Ѓ�_^3�[��]Ë�5���   �J8�E�P�ы�5�����   ��M�Q�҃�_��^[��]��������������U���$SVW3��E��P�M��}܉}��E��  �}��}��O  W�M�Q�U�R���Tr  ���M����wA  ��t��5���   ��U�R�Ѓ�_^3�[��]Ë�5���   �J8�E�P�ы�5�����   ��M�Q�҃�_��^[��]��������������������t��t��t3�ø   ����U���$��5�UVW3���}܉}䋈�   �I,R�E�P�у��U�R�M��E��  �}��}��*N  j�E�P�M�Q���q  �M��@  ��5���   ��M�Q�҃�_^��]� ��U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��M  j�U�R�E�P���q  �M��&@  ��5���   �
�E�P�у�^��]� ��������U���$�EV��M�E�3�Q�M��E�   �E��  �E��E��OM  j�U�R�E�P���p  �M��?  ��5���   �
�E�P�у�^��]� ��������U�조5�H���   ]��������������U�조5�H���   ]�������������̡�5�H���   �⡰5�H���   ��U�조5�H���   V�u�R�Ѓ��    ^]�����������U�조5�H���   ]��������������U�조5�HL�QV�ҋ���u^]á�5�H�U�ER�UP���  RV�Ѓ���u��5�Q@�BV�Ѓ�3���^]����������U�조5�H�U�E���  R�U�� P�ERP�у�]������U�조5�H���   ]��������������U�조5�H�U �ER�UP�ER�UP�ER�UP���   R�Ѓ�]������������̡�5�PL�BLQ�Ѓ���������������̡�5�PL�BPQ�Ѓ����������������U�조5�PL�EP�EPQ�JT�у�]� U�조5�PL�EPQ��  �у�]� �U�조5�PL�EPQ���   �у�]� ̡�5�PL�BXQ�Ѓ����������������U�조5�PL�EP�EP�EPQ�J\�у�]� ������������U���4��5SV��HL�QW�ҋ�3ۉ}�;��x  �M��q  ��5�E�EԋE�]Љ]؉]܉]�]��}̋Q�R0Ph]  �M��ҡ�5���   �BSSW���Ѕ���   ��5�QL�BW�Ћ���;���   ��    ��5���   �B(���ЍM�Qh�   ���u��z��������   �M�;���   ��5���   ���   S��;�tm��5���   �ȋB<V�Ћ�5���   ���   �E�P�у�;�t��5�B@�HV�у���;��\����}��M���,���M��  ��_^[��]� �}���5�B@�HW�ы�5���   ���   �M�Q�҃��M��,���M��a  _^3�[��]� �����̡�5�PL�B`Q�Ѓ���������������̡�5�PL�BdQ�Ѓ����������������U�조5�PL�EPQ�Jh�у�]� ���̡�5�PL��D  Q�Ѓ������������̡�5�PL�BlQ�Ѓ����������������U�조5�PL�EPQ���   �у�]� �U��M��]�����U��M��U�@R��]��������������U��U�M��@R�UR��]����������U��U�M��@R�UR�UR�UR��]��U��U$�EV�Eh�*h�*hp*h`*R�Q�U R�UR�UR�U���A�$�5�5�vLRP���   Q�Ѓ�4^]�  ������̡�5�PL���   Q�Ѓ�������������U�조5�PL�EP�EP�EPQ��   �у�]� ���������U�조5�PL��H  ]�������������̡�5�PL��L  ��U�조5�PL��P  ]��������������U�조5�PL��T  ]��������������U�조5�PL�EP�EP�EP�EP�EPQ���   �у�]� �U�조5�PL�EP�EP�EPQ���   �у�]� ���������U�조5�PL�EP�EP�EP�EPQ��   �у�]� �����U�조5�HL���   ]��������������U�조5�HL���   ]��������������U�조5�HL���   ]�������������̡�5�HL��  �⡰5�HL��@  ��h�5Ph^� ��  ���������������U��Vh�5j\h^� ���  ����t�@\��t
�MQV�Ѓ�^]� ������������U��� ��5V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��5�QLjP���   ���ЋM��U�Rh=���M�}��c������5���   ���   �U�R�Ѓ��M��u��,(����_^��]Ë�5���   ���   �E�P�у��M��u���'��_�   ^��]����U��� ��5V3��u��u�u�u�u��u��u􋈈   ���   W�ҋ}�E�;�t`;�t\��5�QLjP���   ���ЋM��U�Rh<���M�}��������5���   ���   �U�R�Ѓ��M��u��\'����_^��]Ë�5���   ���   �E�P�у��M��u��.'��_�   ^��]���̡�5V�񋈈   ���   V�҃��    ^��������������̸   � ��������� ������������̃��� ����������� �������������U�조5�H�QV�uV�҃���^]� ̸   � ��������3�� ����������̸   @� ��������3��  ����������̸   � ��������U��W�}��u3�_]� ��U�@@VR�Ћ���u^_]� ��5�Q0�F�M���   PQW�ҋF��^_]� U�조5�H0�U�AR�Ѓ���t
��ȋj��]� �������3�� ��������������������������̸   � ��������3�� �����������3�� �����������U��E� ����]� �������������̸   � ��������U��E� ����]� ��������������3�� �����������U�조5�H���  ]��������������U�조5�H���  ]��������������U�조5�P�EP�EP�EP�EPQ���   �у�]� �����U�조5�E�P�EP�E���\$�E�$PQ���   �у�]� �������������U�조5�P�EP�EP�EPQ���   �у�]� ��������̡�5�P���   Q�Ѓ�������������U�조5�P�EP�EP�EPQ���   �у�]� ���������U�조5�P�EP�EPQ���   �у�]� �������������U�조5�H�U�ApR�Ѓ�]� �����U�조5�P�EP�EPQ���  �у�]� �������������U�조5�P�EP�EPQ���  �у�]� �������������U�조5�P�EP�EPQ���  �у�]� �������������U�조5�P�EP�EPQ���  �у�]� �������������U����   V�u��u3�^��]�Wh�   ��0���j P脨  ��R���E�P���ҡ�5�P�B<�M��Ћ}��t0j �M�QW�a#������u��5�B�P�M�Q�҃�_3�^��]ËE�M�Uh�   ��p�����0���P��t����MQWj	��P�����0���ǅ4������E� 7�E� 7�E����E����E�7�E�p��E�@7ǅx�����ǅ|����6�E����E�`7�E�P��E���E�p7�E��6�E����E�07�E�P7�E����EĀ7�	����5���B�P�M�Q�҃�_��^��]����������U���   SV�u(3ۉ]���u��5�H�A�UR�Ѓ�^3�[��]Ë�5�Q�B<W�M3��Ѕ��N  ��B  �E�����   �MQ�M��  ��5�B�P�M�Q�ҡ�5�H�AWj��U�h<�R�Ѓ��M�Q�M��{  �u�Wj��U�R�E�P��\���Q�_?�>   ��P��x���R�n  ��P�E�P�a  ��P����C  �E���t�E� �� t�M�����  ��t��x�������  ��t��\�������s  ��t�M̃���c  ��t��5�Q�J�E�P����у���t�M��9  �}� t"�U(�E$�M�R�UP�EQ�MRPQ����������U�R�A  ����E$�M�UVP�Ej QRP�����������5�Q�J�EP�у���_^[��]���������U��E�M�UP�EQ�Mj RPQ������]�������������̋�`L����������̋�`����������̋�` ����������̋�`0����������̋�`$����������̋�`T����������̋�`����������̋�`����������̋�`8����������̋�`H����������̋�`����������̡�5�P�BVj j����Ћ�^���������U�조5�P�E�RVj P���ҋ�^]� U�조5�P�E�RVPj����ҋ�^]� ��5�P�B�����U�조5�P���   Vj ��Mj V�Ћ�^]� �����������U�조5�P�EPQ�J�у�]� ����U�조5�P�EPQ�J�у����@]� ���������������U�조5�P�E�RtP�ҋ�5���   P�BX�Ѓ�]� ���U�조5�P�E�Rlh#  P�EP��]� ���������������U�조5�P�E�RlhF  P�EP��]� ���������������U�조5�P�E�RtP�ҋ�5���   �M�R`QP�҃�]� ���������������U�조5�P���   ]��������������U�조5�P�E���   P�҅�u]� ��5���   P�B�Ѓ�]� ��������U��E�M�UP��P�EjP�C	����]��������������̸   �����������U��V�u��t���u6�EjP�D	������u3�^]Ë��1
����t���t��U3�;P��I#�^]�������U��� �E�M���  �ȉESHV�u��W�}��A�Q����H։E��B��E���؉M�E��U���I �M��~�U�U�I)}�M��4�E��}���t�u+��\�P@�M���u�EH�E����   )}��u��	;]��u��s���u�]�;]}�M��>P�E�V�Ѕ�y�u�C�]�M��E��VP�҅��d����F��}��t�M�+���I ��P@�M��T�u�]��;]~��/���_^[��]� ������U���(W�}�����E�E�M���/  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��
�U���$    ��~�M�M�J)}��U��G�M�E��M��t'�M�+����$    ��pf�\���M�f�f�4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��H����}�F���t!�M�+ȍI �Pf���Of�f�T�u�]��}�;E�~����	���^[_��]� ����������U���(W�}�����E�E�M���  �ЉEH����B�J���SV�uƃ��ΉE��A��E����؉U��E܉M��	�U���    ��~�M�M�J)}��U��9�M�E��M��t�M�+ȋ\�p���M��4u�EH�E����   )}��u�;E��؉u�s���u�]�;]}�M��>P�E؋V�Ѕ�y�u�C�]��M��E�VP�҅��W����}�F���t�M�+Ȑ��P��O��T�u�]��}�;E~��"���^[_��]� ��U��EP�u�E�UPR����]� 3҅��E�����UPRt	�+���]� �����]� ��������������U����ESV��W�]���t6�u��t/�}��t(�} t"�VP��Ѕ���   xO�E�   �}��}_^3�[��]� �}}���E������uu��VP�҅�tyO�}�G�}��E9E�~�_^3�[��]� ��~3�E���]��]�E����E�M���؋ESPO�҅�u����_��^[��]� �������U����ESV��W�]����  �u����   �}����   �} ��   �VP��Ѕ���   y�M_^�    3�[��]� �O�3��E�   �M��} ����   �EG�8_^3�[��]� �d$ �M�U���<�M������uuVQ���҅�ty�O��M��W�U��M9M�~�뤅�~1�E���]��]�E��E�M���؋ESPO�҅�u����_��^[��]� �M�9_^3�[��]� �U_^�����3�[��]� ������������̡�5V��H�QV�ҡ�5�H$�QDV�҃���^�����������U�조5V��H�QV�ҡ�5�H$�QDV�ҡ�5�U�H$�AdRV�Ѓ���^]� ��U�조5V��H�QV�ҡ�5�H$�QDV�ҡ�5�U�H$�ARV�Ѓ���^]� ��U�조5V��H�QV�ҡ�5�H$�QDV�ҡ�5�H$�U�ALVR�Ѓ���^]� �̡�5V��H$�QHV�ҡ�5�H�QV�҃�^�������������U�조5�P$�EPQ�JL�у�]� ����U�조5�P$�R]�����������������U�조5�P$�Rl]����������������̡�5�P$�Bp����̡�5�P$�BQ�Ѓ����������������U�조5�P$��VWQ�J�E�P�ы�5�u���B�HV�ы�5�B�HVW�ы�5�B�P�M�Q�҃�_��^��]� ���U�조5�P$�EPQ�J�у�]� ����U�조5�P$��VWQ�J �E�P�ы�5�u���B�HV�ы�5�B$�HDV�ы�5�B$�HLVW�ы�5�B$�PH�M�Q�ҡ�5�H�A�U�R�Ѓ� _��^��]� ���U�조5�P$��VWQ�J$�E�P�ы�5�u���B�HV�ы�5�B$�HDV�ы�5�B$�HLVW�ы�5�B$�PH�M�Q�ҡ�5�H�A�U�R�Ѓ� _��^��]� ���U���,VW�E�P�o�����5�Q$�JP�E�P�ы�5�u���B�HV�ы�5�B�HVW�ы�5�B�P�M�Q�ҡ�5�H$�AH�U�R�Ћ�5�Q�J�E�P�у� _��^��]� �����̡�5�P$�B(Q��Yá�5�P$�BhQ��Y�U�조5�P$�EPQ�J,�у�]� ����U�조5�P$�EPQ�J0�у�]� ����U�조5�P$�EPQ�J4�у�]� ����U�조5�P$�EPQ�J8�у�]� ����U�조5�UV��H$�ALVR�Ѓ���^]� ��������������U�조5�H�QV�uV�ҡ�5�H$�QDV�ҡ�5�H$�U�ALVR�Ћ�5�E�Q$�J@PV�у���^]�U�조5�UV��H$�A@RV�Ѓ���^]� ��������������U�조5�P$�EPQ�J<�у�]� ����U�조5�P$�EPQ�J<�у����@]� ���������������U�조5�P$�EP�EPQ�JP�у�]� U�조5�P$�EPQ�JT�у�]� ���̡�5�H$�QX�����U�조5�H$�A\]�����������������U�조5�P$�EP�EP�EPQ�J`�у�]� �����������̡�5�H(�������U�조5�H(�AV�u�R�Ѓ��    ^]��������������U�조5�P(�R]����������������̡�5�P(�B�����U�조5�P(�R]�����������������U�조5�P(�R]�����������������U�조5�P(�R ]�����������������U�조5�P(�E�RjP�EP��]� ��U�조5�P(�E�R$P�EP�EP��]� ��5�P(�B(����̡�5�P(�B,����̡�5�P(�B0�����U�조5�P(�R4]�����������������U�조5�P(�RX]�����������������U�조5�P(�R\]�����������������U�조5�P(�R`]�����������������U�조5�P(�Rd]�����������������U�조5�P(�Rh]�����������������U�조5�P(�Rx]�����������������U�조5�P(�Rl]�����������������U�조5�P(�Rt]�����������������U�조5�P(�Rp]�����������������U�조5�P(�BpVW�}W���Ѕ�t:��5�Q(�Rp�GP���҅�t"��5�P(�Bp��W���Ѕ�t_�   ^]� _3�^]� ��U�조5�P(�BtVW�}W���Ѕ�t:��5�Q(�Rt�GP���҅�t"��5�P(�Bt��W���Ѕ�t_�   ^]� _3�^]� ��U�조5�P(�BpSVW�}W���Ѕ���   ��5�Q(�Rp�GP���҅���   ��5�P(�Rp�GP���҅�tp��5�P(�Bp�_S���Ѕ�tY��5�Q(�Rp�CP���҅�tA��5�P(�Bp��S���Ѕ�t*�OQ��������t��$W��������t_^�   []� _^3�[]� ���U�조5�P(�BtSVW�}W���Ѕ���   ��5�Q(�Rt�GP���҅���   ��5�P(�Rt�GP���҅�tp��5�P(�Bt�_S���Ѕ�tY��5�Q(�Rt�CP���҅�tA��5�P(�Bt��S���Ѕ�t*�O0Q���+�����t��HW��������t_^�   []� _^3�[]� ���U�����5�E�    �E�    �P(�RhV�E�P���҅���   �E���uG��5�H�A�U�R�Ћ�5�Q�E�RP�M�Q�ҡ�5�H�A�U�R�Ѓ��   ^��]� ��5�Qh��h`  P���   �Ћ�5���E��Q(��u�B4j�����3�^��]� �M��Rj QP���҅�u�E�P�������3�^��]� ��5�E��Q�M�j HP�EQ�JP�эU�R�Ĩ�����   ^��]� �����U�조5��V��H�A�U�R�Ѓ��M�Q������^��u��5�B�P�M�Q�҃�3���]� ��5�H$�E�I�U�RP�ы�5�B�P�M�Q�҃��   ��]� �U��Q��5�P(�RX�E�P�҅�u��]� �M3�8E�����   ��]� ���������U�조5�P(�R8]�����������������U�조5�P(�R<]�����������������U�조5�P(�R@]�����������������U�조5�P(�RD]�����������������U�조5�P(�RH]�����������������U�조5�P(�E�R|P�EP��]� ����U�조5�P(�RL]�����������������U�조5�E�P(�BT���$��]� ���U�조5�E�P(�BPQ�$��]� ����̡�5�H(�Q�����U�조5�H(�AV�u�R�Ѓ��    ^]��������������U�조5�P(���   ]��������������U�조5�H(�A]����������������̡�5�H,�Q,����̡�5�P,�B4�����U�조5�H,�A0V�u�R�Ѓ��    ^]�������������̡�5�P,�B8�����U�조5�P,�R<��VW�E�P�ҋu����5�H�QV�ҡ�5�H$�QDV�ҡ�5�H$�QLVW�ҡ�5�H$�AH�U�R�Ћ�5�Q�J�E�P�у�_��^��]� �������U�조5�P,�E�R@��VWP�E�P�ҋu����5�H�QV�ҡ�5�H�QVW�ҡ�5�H�A�U�R�Ѓ�_��^��]� ��̡�5�H,�j j �҃��������������U�조5�P,�EP�EPQ�J�у�]� U�조5�H,�AV�u�R�Ѓ��    ^]�������������̡�5�P,�B����̡�5�P,�B����̡�5�P,�B����̡�5�P,�B ����̡�5�P,�B$����̡�5�P,�B(�����U�조5�P,�R]�����������������U�조5�P,�R��VW�E�P�ҋu����5�H�QV�ҡ�5�H$�QDV�ҡ�5�H$�QLVW�ҡ�5�H$�AH�U�R�Ћ�5�Q�J�E�P�у�_��^��]� �������U�조5�H��D  ]��������������U�조5�H��H  ]��������������U�조5�H��L  ]��������������U�조5�H�I]�����������������U�조5�H�A]�����������������U�조5�H�I]�����������������U�조5�H�A]�����������������U�조5�H�I]�����������������U�조5�H���  ]��������������U�조5�H�A]�����������������U���V�u�E�P���������5�Q$�J�E�P�у���u-��5�B$�PH�M�Q�ҡ�5�H�A�U�R�Ѓ�3�^��]Ë�5�Q�J�E�jP�у���u=�U�R��������u-��5�H$�AH�U�R�Ћ�5�Q�J�E�P�у�3�^��]Ë�5�B�HjV�у���u��5�B�HV�у����I�����5�Q$�JH�E�P�ы�5�B�P�M�Q�҃��   ^��]�����������U�조5�H�A ]�����������������U�조5�H�I(]�����������������U�조5�H��  ]��������������U�조5�H��   ]��������������U�조5�H��  ]��������������U�조5�H��  ]��������������U�조5�H�A$��V�U�WR�Ћ�5�Q�u���BV�Ћ�5�Q$�BDV�Ћ�5�Q$�BLVW�Ћ�5�Q$�JH�E�P�ы�5�B�P�M�Q�҃�_��^��]������U�조5�H���  ��V�U�WR�Ћ�5�Q�u���BV�Ћ�5�Q$�BDV�Ћ�5�Q$�BLVW�Ћ�5�Q$�JH�E�P�ы�5�B�P�M�Q�҃�_��^��]���U�조5�H���  ]��������������U���<��5SVW�E�    ��t�E�P�   �������/��5�Q�J�E�P�   �ы�5�B$�PD�M�Q�҃��}ࡰ5�H�u�QV�ҡ�5�H$�QDV�ҡ�5�H$�QLVW�҃���t)��5�H$�AH�U�R����Ћ�5�Q�J�E�P�у���t&��5�B$�PH�M�Q�ҡ�5�H�A�U�R�Ѓ�_��^[��]���U�조5�H�U���  ��VWR�E�P�ы�5�u���B�HV�ы�5�B$�HDV�ы�5�B$�HLVW�ы�5�B$�PH�M�Q�ҡ�5�H�A�U�R�Ѓ� _��^��]����������������U��V�ujV�a�������^]���������̡�5�H���   ��U�조5�H���   V�uV�҃��    ^]�������������U�조5�P�]�⡰5�P�B����̡�5�P���   ��U�조5�P�R`]�����������������U�조5�P�Rd]�����������������U�조5�P�Rh]�����������������U�조5�P�Rl]�����������������U�조5�P�Rp]�����������������U�조5�P�Rt]�����������������U�조5�P���   ]��������������U�조5�P�Rx]�����������������U�조5�P���   ]��������������U�조5�P�R|]�����������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P�EPQ��  �у�]� �U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U��E��t ��5�R P�B$Q�Ѓ���t	�   ]� 3�]� U�조5�P �E�RLQ�MPQ�҃�]� U��E��u]� ��5�R P�B(Q�Ѓ��   ]� ������U�조5�P�R]�����������������U�조5�P�R]�����������������U�조5�P�R]�����������������U�조5�P�R]�����������������U�조5�P�R]�����������������U�조5�P�R]�����������������U�조5�P�E�R\P�EP��]� ����U�조5�E�P�B ���$��]� ���U�조5�E�P�B$Q�$��]� �����U�조5�E�P�B(���$��]� ���U�조5�P�R,]�����������������U�조5�P�R0]�����������������U�조5�P�R4]�����������������U�조5�P�R8]�����������������U�조5�P�R<]�����������������U�조5�P�R@]�����������������U�조5�P�RD]�����������������U�조5�P�RH]�����������������U�조5�P�RL]�����������������U�조5�P�RP]�����������������U�조5�P���   ]��������������U�조5�P�RT]�����������������U�조5�P�EPQ��  �у�]� �U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P�RX]����������������̡�5�P���   ��U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]��������������U�조5�P���   ]�������������̡�5�P���   ��U�조5�P���   ]�������������̡�5�P���   �ࡰ5�P���   �ࡰ5�P���   ��U�조5�H���   ]��������������U�조5�H��   ]��������������U�조5�H�U�E��VWRP���  �U�R�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�_��^��]������������U�조5�H���  ]��������������U�조5�P(�BPVW�}�Q�]���E�$�Ѕ�tM��5�G�Q(�]�E�BPQ���$�Ѕ�t,��5�G�Q(�]�E�BPQ���$�Ѕ�t_�   ^]� _3�^]� ����U�조5�P(�BTVW�}����$���Ѕ�tE��5�G�Q(�BT�����$�Ѕ�t(��5�G�Q(�BT�����$�Ѕ�t_�   ^]� _3�^]� U��VW�}W��� �����t8�GP���������t)�OQ���������t��$W���������t_�   ^]� _3�^]� ������������U�조5�P(�BTVW�}����$���Ѕ�tr��5�G�Q(�BT�����$�Ѕ�tU��5�G�Q(�BT�����$�Ѕ�t8�OQ���������t)�W0R��������t��HW��������t_�   ^]� _3�^]� ���U�조5�P(�} �R8����P��]� �U�조5�P�BdS�]VW��j ���Ћ�5�Qh���p���   h�  V�Ћ�5���E��u�Q(�B4j�����_^3�[]� �Qj VP�Bh���Ћ�5�Q(�BHV���Ѕ�t ��5�Q(�E�R VP���҅�t�   �3��EP������_��^[]� ������U�조5�U�� V��H$�IWR�E�P�ы�5���B�P�M�Q�ҡ�5�H�A�U�RW�Ћ�5�Q�J�E�P�у��U�R���������5�H�A�U�R�Ѓ�_��^��]� �����������h�5PhD � ������������������U��S�]W�;;�t_3�[]� V�s��u#��u9{u9yuP��uL9QuG^_�   []� �A��u��u9Qu��u'��u#9{�Յ�t��t;�u�C��tċI��t�;�t�^_3�[]� ���������U��EP�d������@]� �����������U��h�5jhD �L�������t
�@��t]��3�]��������Vh�5j\hD ����������t�@\��tV�Ѓ���^�����Vh�5j`hD �����������t�@`��tV�Ѓ�^�������U��Vh�5jdhD ����������t�@d��t
�MQV�Ѓ�^]� ������������U��Vh�5jhhD ���y�������t�@h��t
�MQV�Ѓ�^]� ������������Vh�5jlhD ���<�������t�@l��tV�Ѓ�^�������U��Vh�5h�   hD ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5h�   hD ����������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5jphD ���i�������t�@p��t�MQV�Ѓ�^]� ��5^]� ��U��Vh�5jxhD ���)�������t�@x��t
�MVQ�Ѓ���^]� ����������U��Vh�5jxhD �����������t�@|��t�MVQ�Ѓ�^]� 3�^]� �����U��Vh�5jxhD ����������t�@|��t�MVQ�Ѓ����@^]� �   ^]� ������������̋���������������h�5jhD �O�������t	�@��t��3��������������U��V�u�> t+h�5jhD ��������t�@��tV�Ѓ��    ^]�������U��VW�}���t0h�5jhD ���������t�@��t�MQWV�Ѓ�_^]� _3�^]� ����������U��Vh�5jhD ����������t�@��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�5jhD ���I�������t�@��t�MQV�Ѓ�^]� 3�^]� �����Vh�5j hD ����������t�@ ��tV�Ѓ�^�3�^���Vh�5j$hD �����������t�@$��tV�Ѓ�^�3�^���U��Vh�5j(hD ����������t�@(��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�5j,hD ���Y�������t�@,��t�M�UQRV�Ѓ�^]� 3�^]� �U��Vh�5j(hD ����������t�@0��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������Vh�5j4hD �����������t�@4��tV�Ѓ�^�3�^���U��Vh�5j8hD ����������t"�@8��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���������U��Vh�5j<hD ���I�������t�@<��t
�MQV�Ѓ�^]� ������������Vh�5jDhD ����������t�@D��tV�Ѓ�^�3�^���U��Vh�5jHhD �����������t�M�PHQV�҃�^]� U��Vh�5jLhD ����������u^]� �M�PLQV�҃�^]� �����������U��Vh�5jPhD ���i�������u^]� �M�U�@PQRV�Ѓ�^]� �������Vh�5jThD ���,�������u^Ë@TV�Ѓ�^���������U��Vh�5jXhD �����������t�M�PXQV�҃�^]� U��Vh�5h�   hD �����������u^]� �M�UQ�MR�UQ�MR���   QV�҃�^]� �����U��Vh�5h�   hD ���v�������u^]� �M�UQ�MR���   QV�҃�^]� �������������U��Vh�5h�   hD ���&�������u^]� �M���   QV�҃�^]� �����U��Vh�5h�   hD �����������u^]� �M���   QV�҃�^]� �����U��Vh�5h�   hD ����������u^]� �M���   QV�҃�^]� �����U��Vh�5h�   hD ���f�������t�M�UQ�MR���   QV�҃�^]� ��U���Vh�5h�   hD �%�������u��5�H�u�QV�҃���^��]ËM���   WQ�U�R�Ћ�5�Q�u���BV�Ћ�5�Q�BVW�Ћ�5�Q�J�E�P�у�_��^��]��U��Vh�5h�   hD ����������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   hD ���F�������t���   ��t�MQ����^]� 3�^]� �U��Vh�5h�   hD ����������t���   ��t�MQ����^]� 3�^]� �U��Vh�5h�   hD �����������t���   ��t�MQ����^]� 3�^]� �Vh�5h�   hD ����������t���   ��t��^��3�^����������������U��Vh�5h�   hD ���F�������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������U��Vh�5h�   hD �����������t���   ��t�MQ����^]� ��������U��Vh�5h�   hD ����������t���   ��t�M�UQ�MRQ����^]� 3�^]� ���������Vh�5h�   hD ���i�������t���   ��t��^��3�^����������������VW��3����$    �h�5jphD ��������t�@p��t	VW�Ѓ����5�8 tF��_��^�������U��SW��3�V��    h�5jphD ���������t�@p��t	WS�Ѓ����5�8 tqh�5jphD ��������t�@p��t�MWQ�Ѓ������5h�5jphD �k�������t�@p��t	WS�Ѓ����5V���7�����tG�]����E^��t�8��~=h�5jphD ��������t�@p��t	WS�Ѓ����5�8 u_�   []� _3�[]� ����������U��Vh�5j\hD �����������t3�@\��t,V��h�5jxhD ��������t�@x��t
�MVQ�Ѓ���^]� ��������U��Vh�5j\hD ���i�������t3�@\��t,V��h�5jdhD �G�������t�@d��t
�MQV�Ѓ���^]� ��������U���Vh�5j\hD ����������tG�@\��t@V�ЋEh�5jdhD �E��E�    �E�    ���������t�@d��t
�M�QV�Ѓ���^��]� ���������������U��Vh�5j\hD ����������t\�@\��tUV��h�5jdhD �g�������t�@d��t
�MQV�Ѓ�h�5jhhD �>�������t�@h��t
�URV�Ѓ���^]� ���������������U��Vh�5j\hD �������������   �@\��t~V��h�5jdhD ���������t�@d��t
�MQV�Ѓ�h�5jhhD ��������t�@h��t
�URV�Ѓ�h�5jhhD ��������t�@h��t
�MQV�Ѓ���^]� ��U���Vh�5jthD ���F�������tQ�@t��tJ�MQ�U�VR�Ћu��P���?���h�5j`hD ��������th�@`��ta�M�Q�Ѓ���^��]� h�5j\hD ������u����t4�@\��t-V��h�5jdhD ��������t�@d��th�5V�Ѓ���^��]� ������U���Vh�5h�   hD ���s�������tR���   ��tH�MQ�U�R���ЋuP���k���h�5j`hD �:�������t|�@`��tu�M�Q�Ѓ���^��]� h�5j\hD �E�    �E�    �E�    ������u����t3�@\��t,V��h�5jdhD ���������t�@d��t
�U�RV�Ѓ���^��]� ��������������U�조5���   �BXQ�Ѓ���u]� ��5�Q|�M�RQ�MQP�҃�]� ���U�조5���   �BXQ�Ѓ���u]� ��5�Q|�M�R8Q�MQP�҃�]� ���U��EV��j ���5�Qj j P�B�ЉF����^]� ��̡�5Vj ��H��Aj j R�Ѓ��F^����������������U��V��F��u^]� ��5�Q�MP�EP�Q�JP�у��F�   ^]� ���̡�5�H���   ��U�조5�H���   V�u�R�Ѓ��    ^]����������̡�5�P���   Q�Ѓ�������������U�조5�P�EPQ���   �у�]� ̡�5�H�������U�조5�H�AV�u�R�Ѓ��    ^]��������������U�조5�H�AV�u�R�Ѓ��    ^]��������������U�조5�P��Vh�  Q���   �E�P�ы�5���   �Q8P�ҋ�5���   ��U�R�Ѓ���^��]��������������̡�5�P�BQ�Ѓ����������������U�조5�P�EPQ�J\�у�]� ����U�조5�P�EP�EP�EP�EP�EPQ���   �у�]� �U�조5�P�EP�EP�EP�EPQ�JX�у�]� �������̡�5�P�B Q��Y�U�조5�P�EP�EP�EP�EPQ���   �у�]� �����U�조5�P�EP�EP�EPQ�J�у�]� ������������U�조5�H��   ]��������������U�조5�P�R$]�����������������U�조5�P��x  ]��������������U�조5�P�EP�EP�EP�EPQ�J(�у�]� ��������U�조5�P�E(P�E$P�E P�EP�EP�EP�EP�EP�EPQ�J`�у�(]�$ ����U�조5�P�EP�EP�EP�EPQ�J,�у�]� ��������U�조5V��H�QWV�ҍx���5�H�QV�ҋ�5�Q�M�R4Q�MQ�MQWHPj j V�҃�(_^]� ���������������U�조5�P�E P�EP�EP�EP�EP�EP�EPQ�J4�у� ]� ������������U�조5�P�EP�EPQ�J@�у�]� U�조5�P�EPQ�JD�у�]� ���̡�5�P�BLQ�Ѓ���������������̡�5�P�BLQ�Ѓ���������������̡�5�P�BPQ�Ѓ����������������U�조5�P�EPQ�JT�у�]� ����U�조5�P�EPQ�JT�у�]� ����U�조5�P�EP�EPQ���   �у�]� �������������U�조5�P�E���   ��VP�EPQ�M�Q�ҋu�    �F    ��5���   j P�BV�Ћ�5���   �
�E�P�у� ��^��]� ������̡�5�P�BhQ�Ѓ������������������3��Yp��A`�Ad�Ah�Ax�����A|   ����������������U��E��t�Ap��yd t�Ah]� 3��y|��]� ������̡�5�H�������U�조5�H�AV�u�R�Ѓ��    ^]��������������U�조5�P�E P�EP�EP�EP�EP�EP�EPQ�J�у� ]� ������������U�조5�P�EPQ�J�у�]� ���̡�5�P�BQ��Y�U�조5�P�EP�EPQ�J�у�]� U��VW���d���M�U�x@�EPQR���N���H ���_^]� �U��VW���4���M�U�xD�EPQR������H ���_^]� �V������xH u3�^�W�������΍xH�����H �_^�����U��V�������xL u3�^]� W�������M�U�xL�EPQR������H ���_^]� �������������U��V������xP u���^]� W���o���M�U�xP�EP�EQRP���U���H ���_^]� ��������U��V���5���xT u���^]� W������M�xT�EPQ������H ���_^]� U���S�]VW���t.�M��Ʒ���������xL�E�P�������H ��ҍM�� ����}��tZ��5�H�A�U�R�Ћ�5�Q�J�E�WP�ы�5�B�P�M�Q�҃����y���@@��t��5�QWP�B�Ѓ�_^[��]� ������U��V���E���x` u
� }  ^]� W���-���x`�EP������H ���_^]� ��U��VW������xH�EP�������H ���_^]� ���������U��SVW�������x` u� }  �#������x`�E���P������H ��ҋ���5�H�]�QS�҃�;�A��5�H�QS�҃�;�,���o���M�U�xD�EPQSR���X���H ���_^[]� _^�����[]� ��������������U��V���%���xP u
�����^]� W������M�U�xP�EP�EQ�MR�UPQR�������H ���_^]� ��������������U��V�������xT u
�����^]� W������M�xT�EPQ������H ���_^]� ��������������U��V���u���xX tW���g���xX�EP���Y���H ���_^]� ������������U����MV3��E�PQ�u�u��u�u��u�u��x<  ����t.�E�;�t'��5�J�U�R�U�R�U�R�U�RP�AX�Ѓ�^��]�3�^��]������������̡�5�H��   ��U�조5�H��$  V�u�R�Ѓ��    ^]�����������U�조5�UV��H��(  VR�Ѓ���^]� �����������U�조5�P�EQ��,  P�у�]� �U�조5�P�EQ��,  P�у����@]� �����������̡�5�H��0  �⡰5�H��4  �⡰5�H��p  �⡰5�H��t  ��U��E��t�@�3���5�RP��8  Q�Ѓ�]� �����U�조5�P�EPQ��<  �у�]� �U�조5�P�EP�EP�EPQ��@  �у�]� ���������U�조5�P�EP�EPQ��D  �у�]� �������������U�조5�P�EPQ��H  �у�]� �U�조5�P�E��L  ��VWPQ�M�Q�ҋu����5�H�QV�ҡ�5�H�QVW�ҡ�5�H�A�U�R�Ѓ�_��^��]� ��������������̡�5�P��T  Q�Ѓ�������������U�조5�P�EPQ��l  �у�]� ̡�5�P��P  Q�Ѓ�������������U�조5�P�EPQ��X  �у�]� ̡�5�H��\  ��U�조5�H��`  V�u�R�Ѓ��    ^]�����������U�조5�P�EP�EP�EP�EP�EPQ��d  �у�]� �U�조5�P�EP�EP�EP�EP�EPQ��h  �у�]� �VW���O�4�����3��G �G$�G(�G,�G0�G4�G8�G<�G@�GD�GH�GL�GP�GT�GX�G\�_p��G`�Gd�Gh�Gx�����G|   ��_^����������������V��W�>��t7����	���xP t$S����	��j j �XPj�FP����	���H ���[�    �~` t��5�H�V`�AR�Ѓ��F`    _^������������U��SV��Fx��5�Q��   WV�^dSP�EP�~`W�у��F|����   �> ��   �; ��   �U�~pW�^hSR�t�������u#���h���5�H��0  h�   �҃��E�~P���,����j j jW�^����F|��t��������F|_^[]� �F|_�Fx����^[]� �F|�����    ��5�Q��JP�у��    �F|_^[]� ���V��������3��^p��F`�Fd�Fh�Fx�����F|   ^�������U��QV��~d tg�E;Fxt_�N`W�>�M����;���xP u����(S���(���UR�XP�E�Pj�NQ������H ���[�F|_��u�E�Fx�E��t�    �F`^��]� �M�Fx������t�3�^��]� ���������U��QVW�}����8  ��5�H�QhV�҃�����5u"�H��0  h�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���t�3�9u�~�E���<� t��Q���O6  �EF;u�|�UR�k����_�   ^��]� �������������U��QVW�}�����7  ��5�H�QhV�҃�����5u"�H��0  h�h�  �҃�_3�^��]� �E    �H�U�R�U�EP���   RV�Ѓ���tЋE��t�3�9u�~8��E�<� t'����5�QP�Bh�Ѓ���t�M��R���l5  F;u�|ʍEP�j����_�   ^��]� �������������h�h�   h�5h�   �n������t������3��������V��������N^韶�����������������U��VW�}�7��t�������N�s���V�mm�����    _^]�U���EV���V��������Au��5�H��0  hX�j,�����^��^]� �����U���W������G���U��ȵ������A�  ������A��   ���������AuR������AuKV����U  ����U  �ȅ�u��^����__��]Ëƙ����ʅ�u�u��E�^������__��]���������Au������=����������Au6�����������U������G�����_��������Au�����U����_�
����������-W  �E����U��@���������A{���������__��]�������������__��]����U�����V�E��������At�����������Au������x����@��$�jU  ����x����^�e�����^]� ��������������U����V�E��������u�   �3����]����Az�   �3�3����@�;���W���$����T  ��E���@��$��T  �V����������Au��5�H��0  hX�j�����^����_u������������^]� ���U������EV�ы�������z!��5�؋H��0  hX�j5�����U������$�IT  �]��F�$�;T  �}��$�0T  ��E�$�#T  �^�����&���^��]� ���������������U��M��P]����U��M��P]����U��M��P]����V���̸�F    ��5�HP�h`�VhP�h@��҉F����^����������̃y �̸u��5�PP�A�JP��Y��U��A��u]� ��5�QP�M�Rj Q�MQP�҃�]� ��U��A��t��5�QP�M�RQP�҃�]� ������������U��A��t��5�QP�M�RQP�҃�]� �����������̡�5�HP���   ��U�조5�HP���   ]�������������̡�5�HP�QP�����U�조5�HP�AT]����������������̋��     �@    �V����t)��5�QPP�BL�Ћ�5�QP��J<P�у��    ^�������������U��SV�ً3�W;�t��5�QPP�B<�Ѓ��3�s�}�Eh`�W�C��5�QP�J8hP�h@�P�EP�у��9u~M�I ���z u!���@   ��5�QP���H�RQ�҃���5�HP��A@VR�Ћ�F���A;u|�3�9_^��[]� ��������U��SVW��3�9w~<�]��5�HP��A@VR�Ѓ���t-��5�QPj SjP�B�Ѓ���tF;w|�_^�   []� ��5�QP��JLP�у�_^3�[]� �����������̡�5�PP��JDP�у�������������̡�5�PP��JHP��Y��������������̡�5�PP��JLP��Y���������������U��U�E�@R�URP�I���]� �����3���������������U��V��~ �̸u��5�HP�V�AR�Ѓ��Et	V�^f������^]� ���̋�3ɉH��H�@   �������������U��ыM��tK�E��t��5���   P�B@��]� �E��t��5���   P�BD��]� ��5���   R�PD��]� �����U�조5�P@�Rd]�����������������U�조5�P@�Rh]�����������������U�조5�P@�Rl]�����������������U�조5�P@�Rp]�����������������U�조5���   ���   ]�����������U�조5���   ���   ]����������̡�5�P@�Bt����̡�5�P@�Bx�����U�조5�P@�R|]����������������̡�5�P@���   �ࡰ5���   �Bt��U�조5�P@���   ]�������������̡�5�P@���   ��U�조5�P@���   ]��������������U�조5�P@���   ]��������������U�조5�P@���   ]��������������U�조5�P@���   ]��������������U�조5V��H@�QV�ҋM����t��#�����5�Q@P�BV�Ѓ�^]� �̡�5�PH���   Q�Ѓ�������������U�조5�P@�EPQ�JL�у�]� ���̡�5�P@�BHQ�Ѓ����������������U�조5�P@�EP�EP�EPQ�J�у�]� ������������U�조5�P@�EPQ�J�у�]� ����U�조5�P@�EP�EPQ�J�у�]� U�조5�P@�EPQ�J �у�]� ����U�조5���   �R]��������������U�조5���   �R]��������������U�조5���   �R ]��������������U�조5���   ���   ]�����������U�조5���   ��D  ]�����������U�조5�E���   �E ���   P�E���$P�EP�EP�EP��]� ���������U�조5���   ���   ]����������̡�5���   �B$�ࡰ5�H@�Q0�����U�조5�H@�A4j�URj �Ѓ�]����U�조5�H@�A4j�URh   @�Ѓ�]�U�조5�H@�U�E�I4RPj �у�]�̡�5�H|�������U��V�u���t��5�Q|P�B�Ѓ��    ^]��������̡�5�H|�Q �����U��V�u���t��5�Q|P�B(�Ѓ��    ^]��������̡�5�H@�Q0�����U��V�u���t��5�Q@P�B�Ѓ��    ^]���������U�조5�H@���   ]��������������U��V�u���t��5�Q@P�B�Ѓ��    ^]��������̡�5�PH���   Q�Ѓ�������������U�조5�PH�EPQ��d  �у�]� �U�조5�H �IH]�����������������U��}qF uHV�u��t?��5���   �BDW�}W���Ћ�5�Q@�B,W�Ћ�5�Q�M�Rp��VQ����_^]����������̡�5�P@�BT�����U�조5�P@�RX]�����������������U�조5�P@�R\]����������������̡�5�P@�B`�����U�조5�H��T  ]��������������U�조5�H@�U�A,SVWR�Ћ�5�Q@�J,���EP�ы�5�Z��h��hE  �΋��V���Ph��hE  ���D���P��T  �Ѓ�_^[]����h�5Ph^� � ������������������U��Vh�5jh^� ���ٟ������t�@��t�M�UQRV�Ѓ�^]� 3�^]� �Vh�5jh^� ��蜟������t�@��tV�Ѓ�^�3�^���U��Vh�5jh^� ���i�������t�@��t�M�UQRV�Ѓ�^]� ���^]� U���  Vh�5jh^� ���#�������t/�@��t(�MWQ��x���VR�Ћ��E���b   ���_^��]� �u����a���N`�a�����   �a����   �a����ݞ�  ��^��]� ����U��Vh�5jh^� ��虞������t�@��t�M�UQRV�Ѓ�^]� ��������U��Vh�5jh^� ���Y�������t�@��t�M�UQ�MRQV�Ѓ�^]� ����U��Vh�5j h^� ����������t�@ ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������������U��Vh�5j$h^� ���ɝ������t�@$��t�MQV�Ѓ�^]� 3�^]� �����U��Vh�5j(h^� ��艝������t�@(��t�M�UQ�MR�UQRV�Ѓ�^]� U��QVh�5j,h^� ���H�������t �@,�E���t�E�MPQV�U���^��]� ��^��]� ��������U��Vh�5j0h^� �����������t#�@0��t�E�M�U���$QRV�Ѓ�^]� 3�^]� ��������Vh�5j4h^� ��謜������t�@4��tV�Ѓ�^�3�^���Vh�5j8h^� ���|�������t�@8��tV�Ѓ�^�������U���`Vh�5jDh^� ���F�������t(�@D��t!W�M�VQ�Ћ��E���   ���_^��]� �u����^����^��]� ����U��Vh�5jHh^� ����������t�@H��t
�MQV�Ѓ�^]� ������������U��Vh�5jLh^� ��詛������t�@L��t�MQV�Ѓ�^]� ���^]� ����U��Vh�5jPh^� ���i�������t�@P��t
�MQV�Ѓ�^]� ������������U��Vh�5jTh^� ���)�������t�@T��t
�MQV�Ѓ�^]� ������������U��Vh�5jXh^� ����������t.�@X��t'�M �UQ�MR�UQ�MR�UQ�MRQV�Ѓ� ^]� 3�^]� �������������Vh�5j`h^� ��茚������t�@`��tV�Ѓ�^�3�^���U��Vh�5jdh^� ���Y�������t�@d��t�MQV�Ѓ�^]� 3�^]� �����U���Vh�5jhh^� ����������t1�@h��t*�MQ�U�VR�Ћu��P�������M��������^��]� �u��������^��]� �����������Vh�5jph^� ��謙������t�@p��tV�Ѓ�^Ã��^��Vh�5jlh^� ���|�������t�@l��tV�Ѓ�^Ã��^��Vh�5jth^� ���L�������t�@t��tV�Ѓ�^�3�^���U��Vh�5jxh^� ����������t�@x��t
�MQV�Ѓ�^]� ������������Vh�5j|h^� ���ܘ������t�@|��tV�Ѓ�^�������Vh�5h�   h^� ��詘������t���   ��tV�Ѓ�^�U��Vh�5h�   h^� ���v�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������U��Vh�5h�   h^� ���&�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U���Vh�5h�   h^� ���ӗ������tU���   ��tKW�M�VQ�Ћ�5�u���B�HV�ы�5�B�HVW�ы�5�B�P�M�Q�҃�_��^��]� ��5�H�u�QV�҃���^��]� ����������Vh�5h�   h^� ���9�������t���   ��tV�Ѓ�^Ã��^������������U��Vh�5h�   h^� �����������t���   ��t
�MQV�Ѓ�^]� ������U��Vh�5h�   h^� ��趖������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�5h�   h^� ���f�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������Vh�5h�   h^� ����������t���   ��tV�Ѓ�^�3�^�������������U��Vh�5h�   h^� ���֕������t%���   ��t�M�UQ�MR�UQRV�Ѓ�^]� 3�^]� ���U��Vh�5h�   h^� ��膕������t���   ��t�M�UQRV�Ѓ�^]� ���^]� ����������U��Vh�5h�   h^� ���6�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�5h�   h^� ����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�5h�   h^� ��薔������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�5h�   h^� ���F�������t���   ��t�MQV�Ѓ�^]� ���^]� ��������������Vh�5h�   h^� �����������t���   ��tV�Ѓ�^�3�^�������������Vh�5h�   h^� ��蹓������t���   ��tV�Ѓ�^�3�^�������������Vh�5h�   h^� ���y�������t���   ��tV�Ѓ�^�3�^�������������Vh�5h�   h^� ���9�������t���   ��tV�Ѓ�^�3�^�������������U��Vh�5h�   h^� �����������t!���   ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������Vh�5h�   h^� ��詒������t���   ��tV�Ѓ�^�3�^�������������U���Vh�5h�   h^� ���c�������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�5h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�5h�   h^� ��詑������t���   ��tV�Ѓ�^�3�^�������������U���Vh�5h�   h^� ���c�������tF���   ��t<�MQ�U�VR�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ��U��Vh�5h�   h^� ����������t���   ��t�M�UQRV�Ѓ�^]� ��Vh�5h�   h^� ��詐������t���   ��tV�Ѓ�^�3�^�������������U��Vh�5h�   h^� ���f�������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��QVh�5h�   h^� ����������t#���   �E���t�E�MPQV�U���^��]� ��^��]� ��U��Vh�5h�   h^� ���Ə������t!���   ��t�E�M�U���$QRV�Ѓ�^]� ���������U��Vh�5h�   h^� ���v�������t���   ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�5h�   h^� ���&�������t���   ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5h   h^� ���֎������t��   ��t�MQV�Ѓ�^]� 3�^]� ���������������Vh�5h  h^� ��艎������t��  ��tV�Ѓ�^�3�^�������������U���Vh�5h  h^� ���C�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�5h  h^� ���Í������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U���Vh�5h  h^� ���C�������tB��  ��t8�M�VQ�ЋM���P�Q�P�Q�P�Q�P�@���Q�A��^��]� ��E�P^�P���]� ������U��Vh�5h  h^� ���ƌ������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�5h  h^� ��膌������t��  ��t
�MQV�Ѓ�^]� ������U��Vh�5h  h^� ���F�������t��  ��t
�MQV�Ѓ�^]� ������Vh�5h   h^� ���	�������t��   ��tV�Ѓ�^�3�^�������������U��Vh�5h$  h^� ���Ƌ������t��$  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5h(  h^� ���v�������t!��(  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��Vh�5h,  h^� ���&�������t��,  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�5h0  h^� ���ي������t��0  ��tV�Ѓ�^�3�^�������������U��Vh�5h4  h^� ��薊������t��4  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5h8  h^� ���F�������t��8  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�5h<  h^� �����������t��<  ��t�M�UQ�MRQV�Ѓ�^]� ��������������U��Vh�5h@  h^� ��覉������t��@  ��t�M�UQ�MRQV�Ѓ�^]� ��������������Vh�5hD  h^� ���Y�������t��D  ��tV�Ѓ�^�3�^�������������U��Vh�5hH  h^� ����������t��H  ��t�MQV�Ѓ�^]� 3�^]� ���������������U��Vh�5hL  h^� ���ƈ������t��L  ��t�M�UQRV�Ѓ�^]� 3�^]� �����������U��Vh�5hP  h^� ���v�������t!��P  ��t�M�UQ�MRQV�Ѓ�^]� 3�^]� �������U��QVh�5hT  h^� ���%�������t'��T  �E���t�E�M�UPQRV�U���^��]� ��^��]� ��������������U��Vh�5hX  h^� ���Ƈ������t%��X  ��t�E�M�U���$Q�MRQV�Ѓ�^]� �����U��Vh�5j<h^� ���y�������t�@<��t�M�UQRV�Ѓ�^]� ��������U��Vh�5j@h^� ���9�������t�@@��t�MQV�Ѓ�^]� 3�^]� �����h�5Ph�� � ������������������h�5jh�� �߆������uË@����U��V�u�> t/h�5jh�� 賆������t��U�M�@R�Ѓ��    ^]���U��Vh�5jh�� ���y�������t �@��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jh�� ���)�������t�@��t�M�UQR����^]� ����������U��Vh�5jh�� ����������t�@��t�M�UQR����^]� ����������U��Vh�5jh�� ��詅������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�5j h�� ���Y�������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�5j$h�� ���	�������t �@$��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5j(h�� ��蹄������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5j,h�� ���i�������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  �����������U��Vh�5j0h�� ���	�������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� �������U��Vh�5j4h�� ��蹃������t5�@4��t.�M(�E �UQ�M���$R�UQ�MR�UQ�MRQ����^]�$ 3�^]�$ ������U��QVh�5j8h�� ���X�������t�@8�E���t�E�MPQ���U�^��]� ��^��]� ����������U��Vh�5j<h�� ���	�������t�@<��t�M�UQR����^]� ����������U��Vh�5j@h�� ���ɂ������t�@@��t�M�UQR����^]� 3�^]� ���U��Vh�5jHh�� ��艂������t�@H��t�M�UQR����^]� 3�^]� ���U��Vh�5jDh�� ���I�������t�@D��t�M�UQR����^]� 3�^]� ���U��QVh�5jLh�� ����������t#�@L�E���t�E�EP�����$�U�^��]� ��^��]� �����U��Vh�5jPh�� ��蹁������t�@P��t�M�UQR����^]� 3�^]� ���U��Vh�5jTh�� ���y�������t �@T��t�M�UQ�MR�UQR����^]� 3�^]� �����������U��Vh�5jXh�� ���)�������t(�@X��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��Vh�5j\h�� ���ـ������t(�@\��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ���U��V��~ Wu h�5jh�� 肀������t�@�ЉF�~��t6h�5jh�� �[�������t�@��t�M�UVQ�MRQ����_^]� _3�^]� ��������������U��V��W�~��t+h�5jh�� ��������t�@��t�M�UQR���Ѓ~ t1h�5jh�� ��������t�N�U�M�@R�Ѓ��F    _^]� ����������U��V��~ u h�5jh�� �������t�@�ЉF�v��t+h�5jh�� �\������t�@��t�M�UQR����^]� �������������U��V�q��t@h�5jh�� �������t(�@��t!�M�UQ�MR�UQ�MR�UQR����^]� 3�^]� ��������������U��V�q��t<h�5j h�� �~������t$�@ ��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��SV��~ Wu h�5jh�� �a~������t�@�ЉF�}�]�M�UWSQR���  ��t;�v��t4h�5j$h�� �~������t�@$��t�M�UWSQR����_^[]� _^3�[]� ���U��V�q��t8h�5j(h�� ��}������t �@(��t�M�UQ�MR�UQR����^]� 3�^]� ������U��V�q��tHh�5j,h�� �}������t0�@,��t)�M$�E�UQ�M���\$�E�$R�UQR����^]�  3�^]�  ������U��V�q��t<h�5j0h�� �$}������t$�@0��t�M�UQ�MR�UQ�MRQ����^]� 3�^]� ��U��EHu�E�M��5��5�   ]� �������������U��EHV����   �$�4��   ^]á�5@��5��uT�EP�|����=�.  }�����^]Ëu��t�h�jmh�5j�;������t ���݂����5��tV���,����   ^]���5    �   ^]ËM�UQR�eX���������H^]�^]��W����5u.�3X��认����5��t���]���V�W:������5    �   ^]Ã��^]�P���H�.�ν����h�5Ph�f �{�����������������U��h�5jh�f �l{������t
�@��t]�����]�������U��Vh�5jh�f �;{��������tC�~ t=�E8�M4�U0P�E,Q�M(RPQ���U��R�J����E�NP�у�4�M���t�����^]ÍM�g������^]��U��h�5jh�f ��z������t
�@��t]��3�]��������U��h�5jh�f �z������t�x t�P]��3�]������V��FW��u�~��N�<��u�< ��u_3�^á�5�H�F��  h0�j8��    RP�у���tщ~�F_�   ^���U��V��F;Fu������u^]� �N�V�E���   F^]� �����������U��S�]V��F;�~ ��x�F�M��^�   []� ^3�[]� }jW�F9FuK��u�~��N�<��u�< ��tA��5�B�V��  h0�j8��    QR�Ѓ���t�F�~�N�V��    �F9^|�_�F;Fu���������u����N�V�E���   F^[]� ��U��V��FW�};�~����y3�;Fu�m�����u_^]� �F;�~�N�T����H�;��F�M���F_�   ^]� ����U��E��x2�Q;�}+J�Q;�}V��    �Q�t���@�2;A|�^�   ]� 3�]� ��������������U��Q3�V��~�I�u91t@��;�|���^]� ���������V��W�~W�c3��3����_�F�F^�����A    ��������̋Q�B���x;�}�QV�4���tP�1�����^�3�����������̍Q3��Q�Q�A�Q�A������������W���O�G;�t#��tV�q��t�~ u3���j�ҋ΅�u�^�G�G�G�G    �G�G    _�����U��A��3�V;�t��t�M��B;�t�@��t
�x t��u�3�^]� ����������U��Q�E�P�Q�P�Q�B�A]� �U��E�Q�P�Q�P�Q�B�A]� ̋Q��3�;�t�ʅ�t�I@��t
�y t��u�������������U��E�P�Q�H�A�@�H]� ����U��E�P�Q�H�A�A�H]� ���̋Q��t!�A��t�B�A�Q�P�A    �A    ��������V��W�~W����m1��3����_�F�F^��������������U���SV�uW���^S�}��61��3���F�F�O�N�W���V�E9G~|��I �O���F�U�9FuL��u�~��~��t���< ��tY��5�H���  h0�j8��    RP�у���t0�~�}���V��M����E�F@�E;G|�_^�   [��]� _^3�[��]� U��V�u��x'�A;�} �U��x;�};�t�A��W�<��<���_^]� ���������U��EV�u;�}N��x,�Q;�}%��x!;�};�t�QW�<�P������tVW����_^]� ������������U��V�q3�W��~�Q�}9:t@��;�|����Ѕ�x);�}%N�q;�}�A�t���B�0;Q|�_�   ^]� _3�^]� ������U����E�Qj�E��ARP�M��E����Kx����]� �����U����Q�Ej�E��A�MRPQ�M��E����gx����]� ̋A��;�t?W3�;�t7V�H;�t	9yt���3��P;�t;�t�J�H�P�Q�x�x��;�u�^_������̋Q�,���t!�A��t�B�A�Q�P�A    �A    �̋�� ���@,��HV3��q�q�P�r�r�,��p�p�p�P�H^������V������r����F3��F,�;�t�N;�t�H�F�N�H�V�V�F�F,�;�t�N;�t�H�F�N�H�V�V^�U��E�UP�AR�Ѓ�]� ���������U��V��N3��,�;�t�F;�t�A�F�N�H�V�V�Et	V��0������^]� ������������U��V��W�~W����-��3����E��F�Ft	V�0����_��^]� ������U��V��������Et	V�0������^]� ���������������U�조5�PH�EPQ���  �у�]� �U�조5�P�B4VW�}j��h�  ���ЋMWQ���g��_^]� ��������������U��V���PXW�ҋ}P���ן�����Et�_�   ^]� �M�UPWQR���h��_^]� �����������U��S�]VW��j ��謝���8�  �}uI�~ uC��5�P���   j h�  ���Ѕ�u��5�QP���   h�  ���Ѕ�t	_^3�[]� �M�U�EQ�MRPSWQ���g��_^[]� ��������U��EP�A    ��d����]� �����̸   �A� ������A   � ������U���@S�]VW����`��u�G   �y  ����   �M3�V躜���8�  u4��[��P�w�dd����5�P�M�B4��jh�  ��_^�C�[��]� �MV�u����8�  u�E�M��RPQ����_^�   [��]� �MV�E����8�  t�MV�4����8��  ��5�P�M�B4jh�  �Љw�  ����  �E�H��BXj	��P����3��؃��u�;�t��5�QH���  VS�Ѓ��E��M�;O�b  9w�Y  ��5�B�M���   Vh�  �҅�u!��5�P�M���   Vh�  �Ѕ��  ��5�Q�M�B4Vh�  ��;�t
V���������E��G��5���   ���   �Ћ]�E�;���   ;���   S�b���M���jQ�ˉu��uĉuȉủuЉu؉u���G���U�E��ˉu��u�u�U�E��]��E�   ��V����tHtHt�u���E�   ��E�   ��E�   �ns���M�;�t�"[����BX�M�Q����P�?t���M܃�;�t� [���M������M������M���b���]�U�E�MRSPQ����d��_^[��]� ��5���   ���   �E�P�у�_^�   [��]� �  ��U��V�u����  �����^]� ��U����E�E�EP�M��  h��E�P�E�����  ̋�U��V�u���t  �����^]� ��U����E�E�EP�M��   h��E�P�E����  ̋�U��V�u���'  �����^]� ��U��V����   �EtV�:+��Y��^]� �A��u�ȹË�U��} W��t-V�u�  �pV��  YY�G��t�uVP�  ���G^_]� ��V��~ t	�v��  Y�f �F ^Ë�U��EV��f ����F �0������^]� ��U��V�uW��;�t�����~ t�v���V�����F�G��_^]� ����{�����U��V������h����EtV�A*��Y��^]� ��U��V�u��f ����F �{�����^]� ��Q���!  YË�U��V��������EtV��)��Y��^]� ��U��E��	Q��	P�^  ��Y�Y@]� ��U��� �EVWjY���}��E��E_�E�^��t� t�E� @��E�P�u��u��u�� ��� �����������������������U��WV�u�M�}�����;�v;���  ���   r�=T tWV����;�^_u�4  ��   u������r)��$����Ǻ   ��r����$����$�����$���������#ъ��F�G�F���G������r���$����I #ъ��F���G������r���$����#ъ���������r���$����I w�d�\�T�L�D�<�4��D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$��������������E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$�������$����I �Ǻ   ��r��+��$� ��$���0�T�|��F#шG��������r�����$���I �F#шG�F���G������r�����$����F#шG�F�G�F���G�������V�������$���I ������������ ���D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$����,�4�D�X��E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_�Ë�U��QS�E���E�d�    �d�    �E�]�m��c���[�� XY�$����U��QQSVWd�5    �u��E���j �u�u��u���  �E�@����M�Ad�=    �]��;d�    _^[�� U���SVW��E�3�PPP�u��u�u�u�u�i  �� �E�_^[�E���]Ë�U��V��u�N3��  j V�v�vj �u�v�u�,  �� ^]Ë�U���8S�}#  u���M�3�@�   �e� �E�>��`#�M�3��E��E�E�E�E�E�E�E �E��e� �e� �e� �e�m�d�    �E؍E�d�    �E�   �E�E̋E�E��,!  ���   �EԍE�P�E�0�U�YY�e� �}� td�    ��]؉d�    �	�E�d�    �E�[�Ë�U��QS��E�H3M�  �E�@��ft�E�@$   3�@�l�jj�E�p�E�p�E�pj �u�E�p�u��  �� �E�x$ u�u�u�����j j j j j �E�Ph#  �������E��]�c�k ��3�@[�Ë�U��QSVW�}�G�w�E����+���u�#  �MN��k�E�9H};H~���u	�M�]�u�} }̋EF�0�E�;_w;�v�^#  ��k�E�_^[�Ë�U��EV�u���  ���   �F�  ���   ��^]Ë�U���  ���   �
�;Mt
�@��u�@]�3�]Ë�U��V�u  �u;��   u�e  �N���   ^]��T  ���   �	�H;�t���x u�^]�"  �N�H�ҋ�U����`#�e� �M�3��M�E��E�E�E@�E�4��M��E�d�    �E�E�d�    �uQ�u�"  �ȋE�d�    ����;`#u����"  �s��#��#i���#���#V���#����#��#���#����#=���#��Ë�U�������} t��.  ��]���̃=T ��   ���\$�D$%�  =�  u�<$f�$f��f���d$uU��.  ��=T t2���\$�D$%�  =�  u�<$f�$f��f���d$u�.  ���$�6  �   ��ÍT$�]6  R��<$tmf�<$t�6  =  �?s-����������������=�5 �~6  �   �p#�{6  w8�D$��%�� D$u'��   ���t���������5  ���� u�|$ u����-P��   �=�5 �6  �   �p#�#5  Z����������̃��$��5  �   ��ÍT$�5  R��<$�D$tQf�<$t�@5  �   �u���=�5 ��5  �   ��#�5  �  �u,��� u%�|$ u���5  �"��� u�|$ u�%   �t����-P��   �=�5 �V5  �   ��#�_4  Z�jh�@  �E��uz�j@  ��u3��8  ��  ��u�o@  ����?  ���T�W?  ��5�9  ��y�s  ���>  ��x �<  ��xj �F7  Y��u��5��   �;  ��3�;�u[9=�5~���5�}�9=|9u��8  9}u�`;  �  ��?  �E������   �   3�9}u�=�#�t��  ��j��uY�  h  j�r5  YY��;�����V�5�#�56���Ѕ�tWV��  YY����N��V�I  Y�������uW�*  Y3�@�?  � jh8�F?  ����]3�@�E��u9�5��   �e� ;�t��u.����tWVS�ЉE�}� ��   WVS�C����E����   WVS�F����E��u$��u WPS�2���Wj S��������tWj S�Ѕ�t��u&WVS�������u!E�}� t����tWVS�ЉE��E������E���E��	PQ�A  YYËe��E�����3��>  Ë�U��}u�A  �u�M�U�����Y]� ��U��S�]���woVW�=�: u��C  j�.B  h�   �4  YY��t���3�@Pj �5�:������u&j^9�@tS�sD  Y��u���D  �0�D  �0��_^�S�RD  Y��C  �    3�[]�����̋T$�L$��ti3��D$��u���   r�=T t�8D  W����r1�ك�t+ш����u������������ʃ���t��t
�����u��D$_ËD$Ë�U��} t-�uj �5�:����uV�DC  ����P��B  Y�^]�������������U��WV�u�M�}�����;�v;���  ���   r�=T tWV����;�^_u�  ��   u������r)��$�0��Ǻ   ��r����$�D��$�@���$����T�����#ъ��F�G�F���G������r���$�0��I #ъ��F���G������r���$�0��#ъ���������r���$�0��I '�������������D��D��D��D��D��D��D���D���D��D��D���D���D���D����    ���$�0���@�H�T�h��E^_�Ð���E^_�Ð���F�G�E^_�ÍI ���F�G�F�G�E^_�Ð�t1��|9���   u$������r����$��������$�|��I �Ǻ   ��r��+��$����$�������,��F#шG��������r�����$����I �F#шG�F���G������r�����$�����F#шG�F�G�F���G�������V�������$����I �����������������D��D��D��D��D��D��D��D��D��D��D��D��D��D���    ���$�������������E^_�Ð�F�G�E^_�ÍI �F�G�F�G�E^_�Ð�F�G�F�G�F�G�E^_���5�@����t��j�=  jj �A  ����@  ��U��QSV�5�W�5T���5T�؉]��֋�;���   ��+��G��ruS�A  �؍GY;�sH�   ;�s���;�rP�u���.  YY��u�C;�r>P�u���.  YY��t/��P�4�� ��T�u�= ��׉��V�ףT�E�3�_^[�Ë�Vjj �T.  YY��V� ��T�T��ujX^Ã& 3�^�jhX�b8  ��.  �e� �u�����Y�E��E������	   �E��~8  ���.  Ë�U���u���������YH]�����������̃=T t-U�������$�,$�Ã=T t���<$Xf��f��t�U��� ������T$�|$�l$�T$�D$��t<���y�$�$��   �������� �T$�� �,�$�$������� �T$�� ��T$�����u��\$�\$������̃=T ��B  ���\$�D$%�  =�  u�<$f�$f��f���d$��B  � �~D$f( �f(�f(�fs�4f~�fTP�f��f�ʩ   uL=�  |}f��=2  f�L$�D$�f.�{$��  ���T$�ԃ��T$�T$�$�?  ���D$��~D$f��f(�f��=�  |!=2  �fT��\�f�L$�D$����f�@�fV@�fT0�f�\$�D$���������������̺`��1C  �`��B  ���������z���Ë�U��UVW��t�}��u�8<  j^�0�}F  ���3�E��u����+���@��tOu��u� �<  j"Y�����3�_^]���������������̋L$��   t$�����tN��   u�    ��$    ��$    �����~Ѓ��3�� �t�A���t2��t$�  � t�   �t�͍A��L$+�ÍA��L$+�ÍA��L$+�ÍA��L$+��jhx�	5  j�G  Y�e� �u�N��t/�6�6�E��t9u,�H�JP����Y�v����Y�f �E������
   ��4  Ë���j��E  Y�����̋T$�L$��   u<�:u.
�t&:au%
�t��:Au
�t:au����
�uҋ�3�Ð��������   t���:u��
�t���   t�f���:u�
�t�:au�
�t����W�ƃ�����   �у���te���    fofoNfoV fo^0ffOfW f_0fof@fonPfov`fo~pfg@foPfw`fp���   ���   Ju���tI������t��    fof�v�Ju��t$����t���v�Iu�ȃ�t	��FGIu�X^_]ú   +�+�Q�ȃ�t	��FGIu���t���v�Hu�Y����j
�$��T3������_�����U��V������L����EtV���Y��^]� ��U��VW�}�G��tG�P�: t?�u�N;�t��QR����YY��t3��$�t�t�E� �t�t�t�t�3�@_^]Ë�U��E� � =RCC�t=MOC�t=csm�u*��  ���    ��  ��  ���    ~�  ���   3�]�jh��2  �}�]��   �s��s�u��|  ���   �e� ;utb���~;w|��  �ƋO�4��u��E�   �|� t�sh  S�O�t���  �e� ��u��+���YËe�e� �}�]�u��u���E������   ;ut�s  �s�1  Ë]�u���  ���    ~��  ���   Ë �8csm�u8�xu2�H�� �t��!�t��"�u�x u�  3�A��  ���3��jh���0  �M��t*�9csm�u"�A��t�@��t�e� P�q������E������1  �3�8E��Ëe��e  ̋�U��M�V�uƃy |�Q�I�42���^]Ë�U��3���;�u
�t  �#  �E��E�9~OS�E�V�E�@�@��p� �M�q�P�GE�P�g�������u
K�������E��E�E�E�;|�^[�E���j����C  �  ���    t��  �e� ��  �M���  �]  �Mj j ���   ������j,h8�/  �ً}�u�]�e� �G��E��v�E�P�J���YY�E��  ���   �E��  ���   �E���
  ���   ��
  �M���   �e� 3�@�E�E��u�uS�uW�������E�e� �o�E������Ëe��
  ��   �u�}�~�   �O��O�^�e� �E�;Fsk��T;�~A;L;�F�L�QVj W�������e� �e� �u�E������E    �   �E���.  ��E�맋}�u�E܉G��u�����Y�
  �Mԉ��   �
  �MЉ��   �>csm�uB�~u<�F= �t=!�t="�u$�}� u�}� t�v����Y��t�uV�*���YY�jh`�.  3҉U�E�H;��X  8Q�O  �H;�u�    ��<  � �u��x�t1�U�3�CS�tA�}�w�A  YY����   SV�A  YY����   �G��M��QP�����YY���   �}�E�p�tH�]A  YY����   SV�LA  YY����   �w�E�pV����������   ���t|��W�9Wu8�A  YY��taSV�A  YY��tT�w��W�E�p�d���YYPV�z������9��@  YY��t)SV��@  YY��t�w�@  Y��t�j X��@�E����  �E������E��3�@Ëe��i  3���,  �jh��,  �E�    �t�]�
�H�U�\�e� �uVP�u�}W�F�����HtHu4j�FP�w����YYP�vS�Q�����FP�w����YYP�vS�7����E������m,  �3�@Ëe���
  ̋�U��} t�uSV�u�V������}  �uuV��u ������7�u�uV�����Gh   �u@�u�F�u�KV�u�������(��tVP����]Ë�U���V�u�>  ���   W�  ���    tG�  ���   �H  9t3�=MOC�t*=RCC�t#�u$�u �u�u�u�uV����������   �}� u�1
  �u�E�P�E�PV�u W�X����M���;M�sg���E�S�x�;7|G;p�B���H�Q��t�z u-�Y��@u%�u$�u�u j �u�u�u�u�����u�E����E��M����E�;M�r�[_^�Ë�U���4�MS�]�CVW�E� =�   �I��I�M����|;�|�m	  �u�csm�9>��  �~� ��)  �F;�t=!�t="��  �~ �  �  ���    ��  �  ���   �u�  ���   jV�E��=  YY��u��  9>u&�~u �F;�t=!�t="�u�~ u��  �=  ���    ��   �+  ���   �   �u3����   ����Y��u\3�9~�G�Lh�#�^�����uF��;7|��  j�u�R���YY�EP�M��E���J���h��E�P�E̸��9����u�csm�9>��  �~��  �F;�t=!�t="���  �}� ��   �E�P�E�P�u��u W�����M���;M���   �x�}�M��G��E�9��   ;O���   ��E�G��E��~r�F�@�X� �E��~#�v�P�u�E���������u�M��9E���M�E��}� ��.�u$�}��u �]��u��E��u�u�uV�u�����u�}���E��E����}�;E��P����}�} t
jV�����YY�}� ��   �%���=!���   �����   V�M���Y����   �H  �C  �>  ���   �3  �}$ �M���   Vu�u��u$�����uj�V�u�u�]������v�g����]�{ v&�} ������u$�u �u�S�u�u�uV������ ��  ���    t�6  _^[�Ë�U��V�u�����������^]� ��U��SVW�  ��   �E�M�csm�����"�u �;�t��&  �t�#�;�r
�@ ��   �Aft#�x ��   �} u}j�P�u�u�������j�x u�#ց�!�rX�x tR99u2�yr,9Yv'�Q�R��t�u$V�u �uP�u�u�uQ�҃� ��u �u�u$P�u�u�uQ������ 3�@_^[]�j � ���(�� ��V�5�#�,�����u�56����V�5�#�0���^á�#���tP�5 6���Ѓ�#���#���tP�4���#��6  jh��%  hк�<��u�F\���f 3�G�~�~pƆ�   CƆK  C�Fh )j�}7  Y�e� �vh�8��E������>   j�\7  Y�}��E�Fl��u�)�Fl�vl�9  Y�E������   �T%  �3�G�uj�E6  Y�j�<6  YË�VW���5�#��������Ћ���uNh  j�  ��YY��t:V�5�#�56���Ѕ�tj V�����YY���N���	V�f���Y3�W�@�_��^Ë�V��������uj�k  Y��^�jh 	�W$  �u����   �F$��tP����Y�F,��tP����Y�F4��tP�����Y�F<��tP�����Y�F@��tP�����Y�FD��tP�����Y�FH��tP�����Y�F\=��tP����Yj��5  Y�e� �~h��tW�D���u�� )tW����Y�E������W   j�5  Y�E�   �~l��t#W��7  Y;=)t��@(t�? uW�z8  Y�E������   V�/���Y�#  � �uj�4  YËuj�z4  YË�U��=�#�tK�} u'V�5�#�5,��օ�t�5�#�5�#���ЉE^j �5�#�56�����u�x�����#���t	j P�0�]Ë�Whк�<�����u	�����3�_�V�5H�h�W��h �W�6��h��W�6��h�W�6�փ=6 �50�� 6t�=6 t�=6 t��u$�,��6�4��6|��56� 6�(���#�����   �56P�օ���   �  �56�5 ����56�6���56�6���5 6�6�֣ 6�_2  ��tc�=�h=��56���У�#���tDh  j�N  ��YY��t0V�5�#�56���Ѕ�tj V����YY���N��3�@��i���3�^_�jh(	�?!  �����@x��t�e� ���3�@Ëe��E������(  �X!  ������@|��t������jhH	��   �5$6����t�e� ���3�@Ëe��E������}����hU�� ��$6�������U���SQ�E���E��EU�u�M�m��?  VW��_^��]�MU���   u�   Q�?  ]Y[�� ��U���(  �07�,7�(7�$7�5 7�=7f�H7f�<7f�7f�7f�%7f�-7��@7�E �47�E�87�E�D7��������6  �87�46�(6	 ��,6   �`#�������d#�������\��x6j��>  Yj �X�h��T��=x6 uj�>  Yh	 ��P�P�L��Ë�U��EV���F ��uc������F�Hl��Hh�N�;)t�P.�Hpu��5  ��F;H-t�F�P.�Hpu�D8  �F�F�@pu�Hp�F�
���@�F��^]� ��U���V�u�M��e����u�P��?  ��e�F�P�v>  ��Yu��P�?  Y��xu���M����   �	��	�F�����F��u�^8M�t�E��`p��Ë�U���V�u�M�������E��u���t���   ��:�t@���u��@��t6���et��Et@���u��H�80t����   �	S�:[uH�
@B���u��}� ^t�E��`p��Ë�U����E�����Az3�@]�3�]Ë�U��QQ�} �u�ut�E�P��>  �M��E��M��H��EP�u?  �E�M����Ë�U��j �u�u�u������]Ë�V����tV����@PV�V������^Ë�U��j �u�d���YY]Ë�U��j �u�����YY]Ë�U���SV�u�M�������3�;�u"�F#  j^�0�-  �}� t�E��`p���^[��9Mv�9M~�E�3���	9Ew	�#  j"��W8Mt�U3�9M��3Ƀ:-����ˋ��6����}�?-��u�-�s�} ~�N�E�����   � � F�3�8E��E��}�u����+�]h �SV�=�������ut�N9Et�E�G�80t/�GHy���F-��d|�jd_�� F��
|�j
_�� F�� F��B_t�90uj�APQ�W������}� t�E��`p�3������3�PPPPP�,  ̋�U���,�`#3ŉE��ESV�uW�}j[S�M�Q�M�Q�p�0�?  ����u��!  ��,  ���m�E��t���u��3Ƀ}�-��+�3Ʌ���+��M�Q�NQP3��}�-��3Ʌ�����Q�=  ����t� ��u�E�j P�u��V�u��������M�_^3�[�����Ë�U��j �u�u�u�u�u������]Ë�U���$VW�u�M��E��  3��E�0   �Y���9}}�}�u;�u#��   j^�0�,+  �}� t�E�`p����  9}v؋E��� 9Ew	�   j"�ȋ}��E�G������  S#�3�;���   ����   �E���u�����j �u�^PSW�$�������t�}� � ��  �M�ap��  �;-u�-F�} �0����$�x�Fje��V�)9  YY���U  �} ���ɀ����p��@ �;  %   �3��t�-F�]������$�x����0�F�O�����  �3���'3��u$�F0�O����� ���u�U���E��  ��F1����F�E9Uu���M܋��   �	�	��O����� �M�w;���   �U��E�   �} ~L�W#U���M�#E���� �\>  f��0����9vËM��m���E�����F�Mf�}� �E�M�}�f�}� |Q�W#U���M�#E���� �	>  f��v1�F����ft��Fu� 0H��;Et���9u��:��	�����@��} ~�uj0V������u�E�8 u���} �4����$�p���W�=  3�%�  #�+E�SY�x;�r	�F+����F-������ڋ��0;�|$��  ;�rSQRP�k<  0�F�U�����;�u��|��drj jdRP�E<  0��U�F����;�u��|��
rj j
RP�<  0��U�F���]�0��F �}� t�E�`p�3�[_^�Ë�U���SVW�u���w�ٍM�N�������u#�  j^�0��'  �}� t�E��`p����   �} v׀} t;uu3��?-���f�0 �?-��u�-�s�G��V�^�C���@PVS�J����0�������} ~QV�^����@PVS�&����E����   � � ������y&�߀} u9}|�}�}������Wj0S��������}� t�E��`p�3�_^[�Ë�U���,�`#3ŉE��EVW�}j^V�M�Q�M�Q�p�0�&:  ����u�k  �0�&  ���lS�]��u�S  �0�&  ���S���;�t3Ƀ}�-����+��u�M�Q�M��QP3��}�-���P�^8  ����t� ��u�E�j VS���N�����[�M�_3�^�Y����Ë�U���,�`#3ŉE��EV�uWj_W�M�Q�M�Q�p�0�e9  ����u�  �8��%  ���   �M��t�S�]�3�K�}�-���<0���u��+ȍE�P�uQW�7  ����t� �W�E�H;������|-;E}(��t
�G��u��G��u�E�j�u���u��������u�E�jP�u���u�u������[�M�_3�^�l����Ë�U��E��et_��EtZ��fu�u �u�u�u�u�'�����]Ã�at��At�u �u�u�u�u�u������0�u �u�u�u�u�u�o�����u �u�u�u�u�u�o�����]Ë�U��j �u�u�u�u�u�u�Z�����]Ë�VW3����#� ����#����(r�_^Ë�Vh   h   3�V�j9  ����t
VVVVV�$  ^�j
�$��T3�����������������U�������$�~$�   ��fD$f% �f�fW�f���fs�,f~����    f������� #�- � =�  ��   �YɁ���  �\��Q�fT׃���� �  fU@�fV�f($�@����X��\��Y��Y��Y����X��^�f��f-���\�fs�?��fs�?�Y�fp�Df5���Y��Y���fW��Y�f\%@��Y��X��Y��\�fp���X��\��\�fD$�D$���-�  ��A�-  fs�&fs�&f��fU��\����Y��X�fV��\��Y����\��Q�%�   ������fT�fs�f��fV�fn�fp� ����  ��Y<�@��Y��Y��Y��\�fTP��X��\��X�f-���\��X�f���^�f��fX�@����Y��Y��Y΃��Y��Y��X�f���Y��X��X�% �  f����fp���X��\��X��X��X�fW�fD$�D$����;  = 8  ��   f�f(5��f�f(��f(%��fY�f(-@���fY�fY�fY����Y�fX�fY��Y�fX�fp��fY�fp���\�fp���\��\��\��\��\��X�fD$�D$���-�;  ����   fW�fT= �f%�f(���Y�f(���\�f(��fp�D�Q�fY�fp�Df��fY�fX�f��fY�����Y�fX�fp�D�Y�fTP�fY�fT�fp�D�\��X��Y��\��\��Y�fp���\��^��fX�fY�fp���X�% �  f��fp���X��X��X��X�fW�fD$�D$����� = � ��   f~�fs� f~�������  �?+���� ��   fT$f~�fs� f~с��������  ��� ��   fW�fW���  f���Y��:   ��fD$�T$�ԃ��T$���T$�$�  fD$����fD$�D$���f������fn�fp� f`�fh�fT�fT��X�fD$�D$���f@�fH��X�fD$�D$���fW��Xƺ�  �J��������������̀zuf��\���������?�f�?f��^���٭^����l��剕l����ݽ`���ƅp��� ���a�����������$�����  ��؃��#�zuf��\���������?�f�?f��^���٭^����l��剕l����ݽ`���ƅp��� �Ɋ�a�����ݽ`����Ɋ�a��������Ŋ�$׊���������$�����
�����  ��؃��#��   ������   ����������������۽b���ۭb�����i���@tƅp����ƅp����d����۽b���ۭb�����i���@t	ƅp����ƅp������۽b���ۭb�����i���@t ��۽b���ۭb�����i���@t	ƅp����ƅp�����������-P���p��� ƅp���
��
�t���������U�����E��E�E��E�E��	U�����E��]��M�E�M�E�M�E�M�PQR�'2  ���E�f�}t�m�����������������������������������ËT$��   ��f�T$�l$é   t�   �����   ËB%  �=  �t�ËB��
  ��D$�B�
�����D$�$�,$��
�    �BËD$%  �=  �tËD$�f�<$t�,$Z�f�$f=tf�� t���f�� t�   �����Z��,$ZÃ��$�D$��%  �����$�D$��%  �t==  �t_f�$f=t*f�� u!���f�� t�   ��t����Z��m���Z��,$Z����������������������   s��������������������������   v����떋�U��VW3��u�:�����Y��u'9L9vV�`����  ;L9v��������uʋ�_^]Ë�U��VW3�j �u�u�_1  ������u'9L9vV�`����  ;L9v��������uË�_^]Ë�U��VW3��u�u�1  ��YY��u,9Et'9L9vV�`����  ;L9v��������u���_^]Ë�U��h���<���th��P�H���t�u��]Ë�U���u�����Y�u�d��j�x  Y�j�  YË�V������V��  V�C  V�  V�3  V�1  V�[�����^Ë�U��V�u3����u���t�у�;ur�^]Ë�U��=� th���3  Y��t
�u��Y�����h(�h�����YY��uTVWhG�z�������Y��;�s���t�Ѓ�;�r�=T _^thT�3  Y��tj jj �T3�]�j hh	�V  j�l  Y�e� 3�@9�9��   �|9�E�x9�} ��   �5T�5��֋؉]Ѕ�th�5T�֋��}ԉ]܉}؃��}�;�rK����9t�;�r>�7�֋���������5T�֋��5T��9]�u9E�t�]܉]ЉE؋��}ԋ]���E�,��}�8�s�E� ��t�ЃE����E�<��}�@�s�E�� ��t�ЃE����E������    �} u)��9   j�  Y�u�����} tj�n  Y��h  Ë�U��j j�u������]�jj j ������Ë�U���  �u�  Yh�   ����̋�U���LV�E�P�x�j@j ^V����YY3�;�u����  ��   � S�5�R;�s6���H��f�@� 
�Hf�@ 
�@!
�H3�H/�5 S��@�P���   ;�r�SWf9M��  �E�;��  ����E�þ   �E�;�|��9�R}k�Sj@j �����YY��tQ��R ��   �;�s1���H���` �`��`3 f�@� 
f�@ 

�@/ ���@΍P�;�r҃�9�R|����R3���~r�E�� ���t\���tW�M��	��tM��uP�t���t=����������4� S�E�� ��E�� �Fh�  �FP�p�����   �F�E�G�E�;�|�3ۋ���5 S����t���t�N��q�F���uj�X�
�C�������P�l������tB��t>W�t���t3%�   �>��u�N@�	��u�Nh�  �FP�p���t,�F�
�N@�����C���h����5�R�h�3�_[^�Ã������VW� S���t6��   ;�s!�p�~� tV�|����@   �N�;�r��7�3����' Y���� T|�_^Ã=T u�""  V�5�5W3���u����   <=tGV�x���Y�t���u�jGW�������YY�=`9��tˋ5�5S�3V�G����>=Y�Xt"jS����YY���t?VSP��������uG���> u��5�5�����%�5 �' � T   3�Y[_^��5`9�^����%`9 �����3�PPPPP�  ̋�U��Q�MS3�V���U�   9Et	�]�E��E��>"u3�9E��"��F�E��<���t��B�U���PF�0/  Y��t��} t
�M��E�F�U�M��t2�}� u��� t��	u���t�B� �e� �> ��   �< t<	uF��N��> ��   �} t	�E�E��3�C3��FA�>\t��>"u&��u�}� t�F�8"u���3�3�9E����E����tI��t�\B���u�U���tU�}� u< tK<	tG��t=��P��t#�K.  Y��t��M�E�F��M��E���(.  Y��tF���UF�V�����t� B�U��M�����E^[��t�  ��Ë�U���S3�VW9Tu�  h  ��9VS��:����T�5p9;�t�E�8u�u��U��E�PSS�}��
����E���=���?sJ�M���sB�����;�r6P�������Y;�t)�U��E�P�WV�}�������E���H�T9�5X93�����_^[�Ë�U���SV�����3�;�u3��wf93t��f90u���f90u�W�=��VVV+�V��@PSVV�E��׉E�;�t8P�;���Y�E�;�t*VV�u�P�u�SVV�ׅ�u�u��w���Y�u�S����E��	S���3�_^[�Ë�V�8��8�W��;�s���t�Ѓ�;�r�_^Ë�V�@��@�W��;�s���t�Ѓ�;�r�_^�j h   j ���3Ʌ�����:����5�:����%�: ��h d�5    �D$�l$�l$+�SVW�`#1E�3�P�e��u��E��E������E��E�d�    ËM�d�    Y__^[��]Q�������̋�U���S�]V�s35`#W��E� �E�   �{���t�N�38�����N�F�38�����E�@f�  �M�U�S��[�E�M���t_�I �[�L��D��E�� �E���t���T  �E���x@G�E��؃��u΀}� t$����t�N�38虻���N�V�3:艻���E�_^[��]��E�    �ɋM�9csm�u)�=�� t h���)  ����t�UjR������M�U��  �E9Xth`#W�Ӌ���  �E�M��H����t�N�38�����N�V�3:�����E��H���  �����9S�O���h`#W���  ������U��V���������2  �N\�U��W9t�����   ;�r���   ;�s9t3���t�P��u3���   ��u�` 3�@��   ����   �MS�^`�N`�H����   j$Y�~\�d9 �����   |� �~d=�  �u	�Fd�   �~=�  �u	�Fd�   �n=�  �u	�Fd�   �^=�  �u	�Fd�   �N=�  �u	�Fd�   �>=�  �u	�Fd�   �.=�  �u	�Fd�   �=� �u	�Fd�   �=� �u�Fd�   �vdj��Y�~d��` Q��Y�^`[���_^]Ë�U��csm�9Eu�uP����YY]�3�]Ë�U����`#�e� �e� SW�N�@��  ��;�t��t	�Уd#�eV�E�P����u�3u����3���3����3��E�P����E�3E�3�;�u�O�@����u��G  ����5`#�։5d#^_[�Ë�U��3��M;��t
@��r�3�]Ë��]Ë�U����  �`#3ŉE�SV�uWV������3�Y�����;��l  j�+  Y���  j��*  Y��u�=6��   ���   �6  hL�h  ��:W�g*  ������   h  ��:VSf��<�����  ��uh�SV�/*  ����t3�PPPPP�]  V��)  @Y��<v*V��)  �ET:��+�j��h�+�SP�)  ����u�h��  VW�w(  ����u������VW�c(  ����u�h  h��W��&  ���^SSSSS�y���j��l���;�tF���tA3��G�����f9Gt@=�  r�S�����P�����P�]�����YP�����PV����M�_^3�[������j�)  Y��tj�)  Y��u�=6uh�   �%���h�   ����YYË�U��E3�;�0$tA��-r�H��wjX]Ë�4$]�D���jY;��#���]��������u��%Ã��������u��%Ã�Ë�U��V������MQ�����Y�������0^]Ë�U��E��@]Ë�U���5�@����t�u��Y��t3�@]�3�]�f��QS������u����t7��$    ffAfA fA0fA@fAPfA`fAp���   HuЅ�t7����t��I f�IHu���t��3���t��IJu���t�AHu�[XË��ۃ�+�3�R�Ӄ�t�AJu���t��IKu�Z�U����7!  ��tj�9!  Y��%tjh  @j�r  ��j�.���̋�U��M��%�U#U��#�ʉ�%]Ë�U��E��@]Ë�U��� �e� Wj3�Y�}��9Eu�B����    �  ����x�MV�u��t��u�����    �b  ����S�����E�;�w�M��u�E��u�E�B   �u�u�P�u��B)  ������t�M�x�E��  ��E�Pj �='  YY��^_�Ë�U���uj �u�u�u�<�����]Ë�U��} u�����    ��  ���]��uj �5�:���]Ë�U���(3��E��E�9�@t�5�R�����V�M��   V;���  ��  ���  �  jZ+���   I��   ����   I��   ����   ItN��	�  �E�   �E�<��M��M�u�]���M��]�Q��]���Y����  ����� "   ��  �E�8��M��M�u�]���M��]�Q��E�   �]���Y�  �E�   �E�8���E�0��M�u��M�]���]���?  �U��E�0��W����E�,��ΉU��E�,��?����E�<��q�����tWItHIt9It ��t���  �E�$���E����E�<��M��u��u����E�<��c����E�   �������E���   �E�   �E���������������   �$�%�E�,���E�0���E�8���E����E���t����E����h����E����\����E�����E�����E����M��u�M����M�]���]�M��]�Q�E�   ��Y��u������ !   �E��^�Ðq$z$�$�$�$�$$$�$$�#�$�$�$��U��QQSV���  V�5�%� :  �EYY�M�ظ�  #�QQ�$f;�uU�8  YY��~-��~��u#�ESQQ�$j�57  ���tVS��9  �EYY�f�ES�����\$�E�$jj�A�8  �]��E�Y�EY������DzVS�9  �E�YY�"�� u��E�S���\$�E�$jj�7  ��^[�����������������U���0���S�ٽ\�����=h. t�w�����8����   [����ݕz������U���U���0���S�ٽ\����=h. t�������8�����8�����S   [��ݕz�����U���0���S�u�u�  ���u�u�  ���ٽ\�����8���������   [�À�8�����=�5 uOݕ0�����p���
�t<�t[<�t?
�t3����r����   f��\���f�� u���f�� tǅr���   �   ٭\�����f��6���f%�f�tf=�tC�f��6���f%�f=�t0�ǅr���   �X������������H�����s4�h��,ǅr���   �P������������@�����v�`�VW��l���C��v�����8���u��u��z������{t�u�}����]���r�����\���SP��l����C��P�j  ��_^�E�����U���0���S�u�u�   ���ٽ\�����8�������������[��U����Sf�Ef��f%�f=�uf���f�]��E�]���E��]��m���E[�Ë�U��E��@]Ë�U���(  �`#3ŉE�S�]W���tS�
  Y������ jL������j P������������������0�����������������������������������������������f������f������f������f������f������f��������������E�M������ǅ0���  �������I��������M�������M�������������\�j ���X�������P�T���u��u���tS�  Y�M�_3�[�v����Ë�Vj� �Vj�������V�P�P�L�^Ë�U���5�@����t]���u�u�u�u�u�����3�PPPPP�������Ë�VW3���@�<��%u���%�8h�  �0���p���tF��$|�3�@_^Ã$��% 3����S�|�V��%W�>��t�~tW��W�ȱ���& Y�����&|ܾ�%_���t	�~uP�Ӄ����&|�^[Ë�U��E�4Ű%���]�jh�	����3�G�}�3�9�:u�M���j����h�   �����YY�u�4��%9t���mj�����Y��;�u�����    3��Pj
�X   Y�]�9u+h�  W�p���uW�����Y�[����    �]���>�W�ܰ��Y�E������	   �E��2����j
�)���YË�U��EV�4Ű%�> uP�#���Y��uj����Y�6���^]�SVW�T$�D$�L$URPQQh�,d�5    �`#3ĉD$d�%    �D$0�X�L$,3�p���t;�T$4���t;�v.�4v�\���H�{ u�h  �C�b  �   �C�t  �d�    ��_^[ËL$�A   �   t3�D$�H3�赩��U�h�p�p�p�>�����]�D$�T$��   �U�L$�)�q�q�q(������]� UVWS��3�3�3�3�3���[_^]Ë���j�  3�3�3�3�3���U��SVWj Rh&-Q�|u  _^[]�U�l$RQ�t$������]� Pd�5    �D$+d$SVW�(��`#3�P�e��u��E������E�d�    Ë�U��3�@�} u3�]Ë�U��SV�58�W�}W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��&t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��_^[]Ë�U��W�}����   SV�5D�W�֋��   ��tP�֋��   ��tP�֋��   ��tP�֋��   ��tP�֍_P�E   �{��&t	���tP�փ{� t
�C��tP�փ��Mu֋��   �   P��^[��_]Ë�U��SV�u���   3�W;�to=�/th���   ;�t^9uZ���   ;�t9uP舭�����   ��5  YY���   ;�t9uP�g������   �n5  YY���   �O������   �D���YY���   ;�tD9u@���   -�   P�#������   ��   +�P�������   +�P�������   ����������   =�&t9��   uP�t1  ���   �ά��YY�~P�E   ���&t�;�t9uP詬��Y9_�t�G;�t9uP蒬��Y���Mu�V胬��Y_^[]Ë�U��W�}��t;�E��t4V�0;�t(W�8�j���Y��tV������> Yu��@(tV�s���Y��^�3�_]�jh�	�J����������P.�Fpt"�~l t�����pl��uj �#���Y���]����j�-���Y�e� �5)��lV�Y���YY�E��E������   �j�&���Y�u��-�  t"��t��tHt3�ø  ø  ø  ø  Ë�VW��h  3��FWP�����3��ȋ��~�~�~����~���� )���F+ο  ��@Ou���  �   ��@Nu�_^Ë�U���  �`#3ŉE�SW������P�v����   ����   3�������@;�r�����ƅ���� ��t0���������;�w+�@P������j R�4������C����u�j �v�������vPW������Pjj �7  3�S�v������WPW������PW�vS��5  ��DS�v������WPW������Ph   �vS�5  ��$3���E������t�L���������t�L ��������  ���  @;�r��R��  ǅ��������3�)�������������  ЍZ ��w
�L�Q ���w�L �Q����  A;�rƋM�_3�[�q�����jh�	�����,������P.�Gpt�l t�wh��uj ����Y��������j����Y�e� �wh�u�;5H-t6��tV�D���u�� )tV�#���Y�H-�Gh�5H-�u�V�8��E������   뎋u�j�\���YË�U���S3�S�M������dB���u�dB   �İ8]�tE�M��ap��<���u�dB   ����ۃ��u�E��@�dB   ��8]�t�E��`p���[�Ë�U��� �`#3ŉE�S�]V�uW�d�����3��};�u������3��  �u�3�9�P-��   �E��0=�   r����  �t  ����  �h  ��P�Ȱ���V  �E�PW������7  h  �CVP�W���3�B���{�s9U���   �}� ��   �u�����   �F����   h  �CVP�����M��k�0�u���`-�u��+�F��t)�>����E���L-D;�FG;�v�}���> uЋu��E����}��u�r�ǉ{�C   �i���j�C�C��T-Zf�1f�0����Ju������������L@;�v����~� �0����C��   �@Iu��C�����C�S��s3��ȋ�����{����95dB�T�������M�_^3�[�h�����jh�	�����M���������}�������_h�u�q����E;C�W  h   �����Y�؅��F  ��   �wh���# S�u����YY�E�����   �u��vh�D���u�Fh= )tP�����Y�^hS�=8����Fp��   �P.��   j����Y�e� �C�tB�C�xB�C�|B3��E��}f�LCf�EhB@��3��E�=  }�L��@+@��3��E�=   }��  ��H,@���5H-�D���u�H-= )tP�B���Y�H-S���E������   �0j����Y��%���u �� )tS����Y�p����    ��e� �E��]���Ã=T uj��V���Y�T   3�����������U��SVWUj j h�7�u��j  ]_^[��]ËL$�A   �   t2�D$�H�3��e���U�h�P(R�P$R�   ��]�D$�T$��   �SVW�D$UPj�h�7d�5    �`#3�P�D$d�    �D$(�X�p���t:�|$,�t;t$,v-�4v���L$�H�|� uh  �D��I   �D��_   뷋L$d�    ��_^[�3�d�    �y�7u�Q�R9Qu�   �SQ�@.�SQ�@.�L$�K�C�kUQPXY]Y[� ��Ã%�R ��U��W�}3�������ك��E���8t3�����_�Ë�U����u�M������E����   ~�E�Pj�u��/  ������   �M�H���}� t�M��ap��Ë�U��=�B u�E�)�A��]�j �u����YY]Ë�U���SV�u�M������]�   ;�sT�M胹�   ~�E�PjS�r/  �M������   �X����t���   ��   �}� t�E��`p����   �E胸�   ~1�]�}�E�P�E%�   P��/  YY��t�Ej�E��]��E� Y������ *   3Ɉ]��E� A�E�j�p�U�jRQ�M�QV�p�E�P�W-  ��$���o������E�t	�M�����}� t�M��ap�^[�Ë�U��=�B u�E�H���w�� ]�j �u�����YY]Ë�U���(�`#3ŉE�SV�uW�u�}�M��?����E�P3�SSSSW�E�P�E�P��9  �E�E�VP�"/  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�Қ���Ë�U���(�`#3ŉE�SV�uW�u�}�M�藾���E�P3�SSSSW�E�P�E�P�)9  �E�E�VP��3  ��(�E�u+��u8]�t�E�`p�jX�/��u8]�t�E�`p�j���E�u��E�u�8]�t�E�`p�3��M�_^3�[�*����Ë�U��MS�YV�u3�;�u����j^�0��������   9Ev�U�;�~��@9Ew�p���j"Y�����W�~�0�ǅ�~���t��C�j0Y�@J���M�  ��x�;5|�� 0H�89t�� �>1u�A�W�3���@PWV�:�����3�_^[]Ë�U��Q�M�AS����% �  V��  #�W�E�A�	���   �%�� �u���t;�t�� <  �(��  �$3�;�u;�u�Ef�M�P��B��<  �U����������U��E����������Ɂ���  ��P��t�M�_^f�H[�Ë�U���0�`#3ŉE��ES�]V�E�W�EP�E�P�"���YY�E�Pj j���uЋ���f���=  �u܉C�E��E��C�E�P�uV虥����$��u�M�_�s^��3�[�C�����3�PPPPP���������������������WVU3�3�D$�}GE�T$���ڃ� �D$�T$�D$�}G�T$���ڃ� �D$�T$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�؋L$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$My���؃� �ʋӋًȋ�Ou���؃� ]^_� ̀�@s�� s����Ë�3Ҁ����3�3��j�m���YË�U��E�M%����#�V�u������t$��tj j �F  YY��x���j^�0�������P�u��t	�gF  ���^F  YY3�^]Ë�S��QQ�����U�k�l$���   �`#3ŉE��C�V�s�HW��x���tRHtCHt4Ht%HtFHHtH��   ǅ|���   �9�   �   ǅ|���   �"ǅ|���   �ǅ|���   �
ǅ|���   Q�~W��|����  ����uI�C��t��t��t�e����M��F����]����M�W�NQP��|�����x���P�E�P�D  ��h��  ��x�����  �>YYt�=h. uV�<  Y��u�6�  Y�M�_3�^膕����]��[Ë�U��M��tj�3�X��;Es������    3�]��MV���uF3����wVj�5�:����u2�=�@ tV�
���Y��uҋE��t�    3���M��t�   ^]Ë�U��} u�u�����Y]�V�u��u�u�����Y3��MW�0��uFV�uj �5�:�̰����u^9�@t@V����Y��t���v�V�{���Y�����    3�_^]���������P����Y������������P����Y����ʋ�U��E��B��B��B��B]Ë�U��E���V9Pt��k�u��;�r�k�M^;�s9Pt3�]��5�B���j h
�-���3��}�}؋]��Kt��jY+�t"+�t+�tY+�uC�������}؅�u����T  ��B��B�U�w\���]���Y�p��Q�Ã�t2��t!Ht�����    �F���빾�B��B���B��B�
��B��B�E�   P���E�3��}���   9E�uj�D���9E�tP�x���Y3��E���t
��t��u�O`�MԉG`��u>�Od�M��Gd�   ��u,����M܋����9M�}�M�k��W\�D�E����ȯ����E������   ��u�wdS�U�Y��]�}؃}� tj �	���Y�S�U�Y��t
��t��u�EԉG`��u�EЉGd3������Ë�U��E��B]�������̋�U��M�MZ  f9t3�]ËA<��8PE  u�3ҹ  f9H��]�����������̋�U��E�H<��ASV�q3�W�D��t�}�H;�r	�X�;�r
B��(;�r�3�_^[]������������̋�U��j�h(
h d�    P��SVW�`#1E�3�P�E�d�    �e��E�    h   �*�������tT�E-   Ph   �P�������t:�@$���Ѓ��E������M�d�    Y_^[��]ËE�3ҁ9  ���Ëe��E�����3��M�d�    Y_^[��]Ë�U����u�M��ô���E�M�U�Tu�} t�M����   �A#E�3���t3�@�}� t�M��ap��Ë�U��jj �uj ������]Ë�U���$�`#3ŉE��ES�E��EVW�E��v����e� �=�B �E�u}hH��а�؅��  �=H�h<�S�ׅ���   �5 �P��h,�S��B��P��h�S��B��P��h��S��B��P�֣�B��th��S��P�֣�B��B�M�5�;�tG9�Bt?P���5�B���֋؅�t,��t(�ׅ�t�M�Qj�M�QjP�Ӆ�t�E�u	�M    �3��B;E�t)P�օ�t"�ЉE��t��B;E�tP�օ�t�u��ЉE��5�B�օ�t�u�u��u��u����3��M�_^3�[�����Ë�U��V�uW��t�}��u����j^�0�������_^]ËM��u3�f��݋�f�: t��Ou��t�+��f�
��f��tOu�3���u�f��5���j"Y���몋�U��US�]VW��u��u9Uu3�_^[]Å�t�}��u�����j^�0�?������݅�u3�f��ЋM��u3�f��ԋ��u��+��f���f��t'Ou��"��+��f���f��tOtKu��u3�f����y���3����u�MjPf�DJ�X�d���f��k���j"Y����j�����U��Ef���f��u�+E��H]Ë�U��V�uW��t�}��u�*���j^�0�o�����_^]ËE��uf��ߋ�+��f���f��tOu�3���u�f������j"Y���뼋�U��M��x��~��u�6]á6�6]������    ��������]Ë�U��E��t���8��  uP����Y]Ë�U��QV�uV�NK  �E�FY��u�b���� 	   �N ����/  �@t�G���� "   ��S3ۨt�^���   �N�����F�F�����F�^�]��  u,�+I  �� ;�t�I  ��@;�u�u�H  Y��uV�fH  Y�F  W��   �F�>�H��N+�I�N;�~WP�u�bG  ���E��M�� �F����y�M���t���t����������� S���#�@ tjSSQ�0?  #����t%�F�M��3�GW�EP�u��F  ���E�9}�t	�N �����E%�   _[^���A@t�y t$�Ix��������QP�v���YY���u	��Ë�U���G@SV����t2� u,�E�+��M������C�>�u�����8*u�ϰ?�����} �^[]Ë�U���x  �`#3ŉE�S�]V�u3�W�u�}������������������������������������������������������������蕮����u+�.����    �r��������� t
�������`p������
  �F@u^V��H  Y��#���t���t�ȃ�������� S����A$u����t���t�ȃ������ S����@$��q���3�;��g����3ɉ��������������������������:
  G������9������'
  �B�<Xw����X����3����x�j��Y������;���	  �$��V��������������������������������������������	  �� tJ��t6��t%HHt���v	  �������j	  �������^	  �������R	  �������   �C	  �������7	  ��*u,���������[�������;��	  �������������	  ������k�
�ʍDЉ�������  ��������  ��*u&���������[�������;���  ��������  ������k�
�ʍDЉ������  ��ItU��htD��lt��w��  ������   �s  �?luG������   �������X  �������L  ������ �@  �<6u�4u�������� �  �������  <3u�2u�������������������  <d��  <i��  <o��  <u��  <x��  <X��  ������������ ������P��P�+  Y��������Yt"������������������G������������������������������i  ��d��  �y  ��S��   ��   ��AtHHtXHHtHH��  �� ǅ����   ������������@�������   ������������9������H  ǅ����   �  ������0  ��   ������   �   ������0  u
������   ���������u������������  �������[���������  ;�u�d.������������ǅ����   �y  ��X��  HHty+��'���HH��  ��������  ������t0�C�Ph   ������P������P��E  ����tǅ����   ��C�������ǅ����   �������������/  ���������;�t;�H;�t4������   � ������t�+���ǅ����   ��  ��������  �`.������P�����Y��  ��p��  ��  ��e��  ��g�4�����itq��nt(��o��  �������ǅ����   ta������   �U�3���������wC  ���:��������� tf������f���������ǅ����   ��  ������@ǅ����
   �������� �  ��  ��S����  u��gucǅ����   �W9�����~�������������   ~=��������]  V�
���������Y��������t���������������
ǅ�����   ��5����������C�������������P��������������������P������������WP�5�#���Ћ���������   t������ u������PW�5�#����YY������gu��u������PW�5�#����YY�?-u������   G������W�
���ǅ����   �������$��s�����HH���������  ǅ����'   �������ǅ����   �p���������Qƅ����0������ǅ����   �L�����   �R������� t��������@t�C���C����C���@t��3҉�������@t��|��s�؃� �ځ�����   ������ �  �ڋ�u3ۃ����� }ǅ����   ���������   9�����~���������u!������u����������������t-�������RPSW�C  ��0���������ڃ�9~������N뽍E�+�F������   ������������tb��t�΀90tW�������������0@�?If90t��;�u�+��������(;�u�`.�������������I�8 t@;�u�+����������������� �~  �������@t2�   t	ƅ����-��t	ƅ����+��tƅ���� ǅ����   ������+�����+������������u'����~!������������� O�m����������t����������������������������v���������Yt(������u��������ϰ0K�����������t��ヽ���� ������tW��~S�������Pj�E�P������PK���i@  ����u#9�����t�������������M������Y��u����������������S�����������Y������ |.������t%��������������ϰ K�n����������t��ヽ���� t���������������� Y���������������t������������3�������������� t
�������`p��������M�_^3�[����Ë��N�L�LJM�M�M�MO3�Ë�U��E�MSVW3��x�E3ۉx�EC�x��t�E	X�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ���t�E�H�E�  ��u��E����3H��1H��E���3H��1H��E����3H��1H��E����3H��1H��E����3H#�1H�  ��t�M�I�t�M�I�t�M�I�t�M�I� t�E	X��   #�t5=   t"=   t;�u)�E��!�E���������E��������E� ���   #�t =   t;�u"�E� ���E�������E�������E�M��3���� 1�E	X 9} �E�}t&�` �E� �E�X�E	X`�E�``���E�XP�4�H �����H �E� �E�X�E	X`�E�H`�����H`��E�XP�c  �EPSj �u� ��M�At�&��At�&��At�&��At�&�Yt�&ߋ��3�+ú����t/HtHtHu(�   � �%����   ���%����   ��!�����+�tHtHu!��#�   �	�#�   �9] t�AP���AP�_^[]Ë�U��j �u�u�u�u�u�u������]Ë�U����ESV3ۋ���C�u��t�]tS�  Y����  �t�Etj�y  Y����x  ����   �E��   j�W  �EY�   #�tT=   t7=   t;�ub��M����h/��{L�H��M�����{,�h/�2��M�����z�h/���M�����z�X/��X/��������   ���   �E��   3��t��W�}���������D��   ��E�PQQ�$�  �M��]�� �����������}�E�����S���]�����Au���3ҋE����f�E����;�}"+��]�t��u���m�]�t�M�   ��m�Hu���t�E����]��E�����_��tj�   Y�e���u��Et�E tj ��  Y���3���^��[�Ë�U��}t~�}������ "   ]������� !   ]Ë�U��E� tj��t3�@]ètj��tjX]������]Ë�U��� 3���p.;Mtd@��|�3��E��t^�E�E�E�E�E�E��EV�u�E�E �E��E$h��  �u(�u��E���  �E�P�S�������uV�,���Y�E�^�Ë�t.�h��  �u(�  �u�����E ���Ë�U��=h. u(�u�E���\$���\$�E�$�uj�/�����$]������h��  �u� !   �\  �EYY]Ë�S��QQ�����U�k�l$���   �`#3ŉE��s �CP�s��������u#�e��P�CP�CP�s�C �sP�E�P�j������s�o������=h. u+��t'�s �C���\$���\$�C�$�sP�q�����$�P�����$��  �s �  �CYY�M�3��dx����]��[Ë�U��QQ�E���]��E��Ë�U��QQ�E�E�M�]��  �����  �f�E��E��Ë�U��3ҁ}  �u
9Uu3�@]Á}  ��u
9UujX]�f�M��  V��f#�^f;�uj���  f;�u�E�� u9Utj��3�]Ë�U���E������������Dz3��   �E3ɩ�  uk�E�� u9Mt]�]��������Au3�@�3���e�E   �t�M�eJ�Et�V���  f!u^;�t	� �  f	E�EQQQ�$��������&Q���EQQ�$������U�����  �����  �E�]Ë�U��Q��}��E��Ë�U��Q�}����E��Ë�U��Q��}��E�M#M��f#E�f����E�m�E��Ë�U��QQ�M��t
�-�/�]���t����-�/�]�������t
�-�/�]����t	�������؛�� t���]����jhH
莹��3�9TtV�E@tH9�/t@�E��U�.�E� � =  �t
=  �t3��3�@Ëe�%�/ �e��U�E�������e��U�n������������V�D$�u(�L$�D$3���؋D$������d$�ȋ��d$��G�ȋ\$�T$�D$���������u�����d$�ȋD$���r;T$wr;D$v	N+D$T$3�+D$T$���؃� �ʋӋًȋ�^� ��U��V�u���c  �v�L{���v�D{���v�<{���v�4{���v�,{���v�${���6�{���v �{���v$�{���v(�{���v,��z���v0��z���v4��z���v��z���v8��z���v<��z����@�v@��z���vD��z���vH�z���vL�z���vP�z���vT�z���vX�z���v\�z���v`�z���vd�z���vh�zz���vl�rz���vp�jz���vt�bz���vx�Zz���v|�Rz����@���   �Dz�����   �9z�����   �.z�����   �#z�����   �z�����   �z�����   �z�����   ��y�����   ��y�����   ��y�����   ��y�����   ��y�����   ��y�����   �y�����   �y�����   �y����@���   �y�����   �y�����   �{y�����   �py�����   �ey�����   �Zy�����   �Oy�����   �Dy�����   �9y�����   �.y�����   �#y�����   �y�����   �y����   �y����  ��x����  ��x����@��  ��x����  ��x����  ��x����  �x����  �x����   �x����$  �x����(  �x����,  �x����0  �{x����4  �px����8  �ex����<  �Zx����@  �Ox����D  �Dx����H  �9x����@��L  �+x����P  � x����T  �x����X  �
x����\  ��w����`  ��w����^]Ë�U��V�u��tY�;�/tP��w��Y�F;�/tP�w��Y�F;�/tP�w��Y�F0;�/tP�w��Y�v4;5�/tV�w��Y^]Ë�U��V�u����   �F;�/tP�cw��Y�F;�/tP�Qw��Y�F;�/tP�?w��Y�F;�/tP�-w��Y�F;�/tP�w��Y�F ;�/tP�	w��Y�F$;�/tP��v��Y�F8;�/tP��v��Y�F<;�/tP��v��Y�F@;�/tP��v��Y�FD;�/tP�v��Y�FH;�/tP�v��Y�vL;5�/tV�v��Y^]Ë�U����`#3ŉE��US3�VW;�~�E��I8t@;�u������+�H;�}@�E�]�9]$u�E� �@�E$�5ذ3�9](SS�u���u��   P�u$�֋��}�;�u3��R  ~Cj�3�X����r7�D?=   w�l"  ��;�t� ��  �P�t��Y;�t	� ��  ���E���]�9]�t�W�u��u�uj�u$�օ���   �5԰SSW�u��u�u�։E�;���   �   �Mt)�E ;���   9E���   P�uW�u��u�u���   �}�;�~Bj�3�X����r6�D?;�w�!  ��;�th���  ���P�t��Y;�t	� ��  �����3�;�t?�u�W�u��u��u�u�օ�t"SS9] uSS��u �u�u�WS�u$����E�W����Y�u��~����E�Y�e�_^[�M�3��}n���Ë�U����u�M��U����u(�E��u$�u �u�u�u�u�uP�������$�}� t�M��ap��Ë�U��QQ�`#3ŉE�S3�VW�]�9]u�E� �@�E�5ذ3�9] SS�u���u��   P�u�֋�;�u3��~<�����w4�D?=   w�p   ��;�t� ��  �P��r��Y;�t	� ��  ���؅�t��?Pj S�<s����WS�u�uj�u�օ�t�uPS�u�ܰ�E�S�Q����E�Y�e�_^[�M�3��Pm���Ë�U����u�M��(����u$�E��u�u�u�u�uP��������}� t�M��ap��Ë�U���S�u�M������]�C=   w�E苀�   �X�u�]�}�E�P�E%�   P�o   YY��t�Ej�E��]��E� Y�
3Ɉ]��E� A�E�j�p�p�E�PQ�E�P�E�jP�6����� ��u8E�t�E��`p�3���E�#E�}� t�M��ap�[�Ë�U����u�M��0����E�M����   �A% �  �}� t�M��ap��Ë�U��j �u����YY]Ë�U���8�`#3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=0O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�0��+0;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�50N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��0�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �0;0��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�003�@�   0�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+0��M���Ɂ�   �ً0]���@u�M̋U�Y��
�� u�M̉�M�_3�[�f���Ë�U���8�`#3ŉE��E�M�M��H
S�ف� �  �MȋH�M��H� ���  ���?  ��W�M�E������u'3�3�9\��u@��|�3��  3��}�j�X�  �e� V�u��}䥥��=(0O�G�������W��  ��]ԉE�yJ���B�t��j3�Y+�@���MЅ��   �E؃�����҅T����|�� u@��|��n�ǙjY#������  �yO���G�e� +�3�B��L���9��}��99}�r"9U����t+�e� �L����z�}�;�r��s�E�   H�U���M�yщM܋MЃ����jY!�E�@;�}
�|��+�3��}� tC�$0��+(0;�}3��}𫫫�	  ;��  +Eԍu�ȍ}𥙃�¥������  ��yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�5(0N�F�������V��  ��E�yJ���BjY+�3�B��\���Mԅ��   ������҅T����|�� u@��|��f�ƙjY#������  �yN���F�e� 3�+�B��L���1�<;�r;�s�E�   �9�M����t�L����r3�;�r��s3�G�1��HyދMԃ����!�E�@��}jY�|��+�3��,0�A���Q����  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�j3�X�S  �,0; 0��   3��}𫫫�M�   �����������  �yJ���B�e� �e� ��������E�    )U��׋]��\���3��#ωMԋ���M�u؉3�u����E��}��u�|Ӌ�j���M�Z+�;�|�1�t����d�� ��Jy�40 03�@�   40�e��������������  �yJ���B�e� �e� ��������E�    )U��֋M��|����#ΉMԋ���M�}؉|���}ԋM����E��}��}�|Ћ�j���M�Z+�;�|�1�t����d�� ��Jy�3�^jY+,0��M���Ɂ�   �ً00]���@u�M̋U�Y��
�� u�M̉�M�_3�[�ka���Ë�U���|�`#3ŉE��E3�V3��E��EFW�E��}��M��u��M��M��M��M��M��M��M�9M$u諪���    ����3��<  �U�U��< t<	t<
t<uB��S�0�B���  �$��{�Hπ�wjYJ�ߋM$�	���   �	:ujY������+tHHt���|  ���jY�E� �  뤃e� jY뛍Hωu���v��M$�	���   �	:uj�<+t"<-t:�t�<C�/  <E~
,d<�!  j�Jj넍Hπ��_����M$�	���   �	:�a���:��s����U��  �u��<9�}�s
�E�*ÈG��E��B:�}�M$�	���   �	:�h���<+t�<-t��k����}� �u��u�u&��M��B:�t��<9Ճ}�s�E�*ÈG�M��B:�}��*Éu�<	�n���j�����J��M��Hπ�wj	��������+t HHt���=���j�����M��jY�Q���j�~����u���B:�t�,1<v�J�&�Hπ�v�:�뿃}  tG����+�J��M�t�HHt��у}� �E����  jX9E�v�}�|�E�O�E��E��}� ��  �Yj
YJ��
�����뾉u�3��<9 k�
���L1Ё�P  	�B:�}���Q  �M��<9�]����B:�}��Q����M��E�O�? t�E�P�u��E�P�  �E�3҃�9U�}��E�9U�uE9U�u+E=P  �!  =�����-  ��2��`�E�;���  }�ع04�E���`9Uu3�f�E�9U���  ��M�3ҋE��}���T���M�;���  k��� �  f9r��}�����M��]��U�3��E��EԉE؉E��C
��3uι�  #�#��� �  ��  ��u���f;��   f;��  ���  f;��	  ��?  f;�w3��EȉE��  3�f;�uA�E����u9u�u9u�u3�f�E���  f;�u!A�C���u9su93u�ủuȉu���  �u��}��E�   �E��U���U���~R�DĉE��C�E��E��U��� �e� �W��4;�r;�s�E�   �}� �w�tf��E��m��M��}� ����E��M��}� ����  f��~7�}܅�x+�u؋E��e����������?���  �u؉E�f���f��M����  f��yB��������E�t�E��E܋}؋U��m�������E������N�}؉E�u�9u�tf�M�� �  f9E�w�Uԁ��� �� � u4�}��u+�e� �}��u�e� ���  f9U�uf�E�A�f�E���E���Eָ�  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�M�f�EċE؉EƋE܉E�f�M��3�f�����e� H%   � ���e� �Ẽ}� �=����E��MċuƋU����/�E�   �3���  �   �3��E�   ��E�   3�3�3�3��}�E�f�f�G
�E��w�W[�M�_3�^��Z���ÍI |u�uvJv�v�v�v4ww�w�w@w��U���t�`#3ŉE��E�U� �  #�S�]�E��A�V#�f�}� W�]��E������E������E����?�E�   t�C-��C �u�}f��u7����   ����   3�f9M�f�����$ �Cf�C0�C 3�@�  f;���   �M3�@f��   �;�u�} t��   @uh���S3�PPPPP�<���3�f9U�t��   �u9Uu-h���;�u"9Uuh���CjP�f������u��C�h���CjP�f������u��C3��k  �ʋ�i�M  �������Ck�M��������3�f�M��ع�2��`�ۉE�f�U�u�}�M���  ��y�04��`�ۉE�����  �E�T�������g  k�M����M�� �  f9r���}ĥ��Eĥ�MƉE�3ɉM��M��M�M��H
��3U��  �� �  �U��U�#�#΍4����  f;���  f;���  ���  f;���  ��?  f;�w3��u�u�u���  3�f;�uG�E����u9u�u9u�u3�f�E��  f;�uG�@���u	9pu90t�!u��u��E�   �M��U�ɉU���~U�L����M��E��E���E�� �V��ȃe� �
;�r;�s�E�   �}� �F�tf��E��m��M��}� ��E����E��M��}� ����  f��~;�E�   �u-�E�M��e��������E�E�������  �E�f���f��M����  f��yB��������E�t�E��M��u�U��m������M������H�u�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�G�f�E���E���E��  f;���   3�3�f9E��E����E�I��   ��� ���M�3�;��}����M�����?  ��  f;���  �]��E�3҉U��U��U�U��U�3�#�#Ё� �  �4
�]���f;��L  f;��C  ���  f;��5  ��?  f;�wK3��E�E��9  f�E�}�f�E��E�E�E��E�f�}��Z���3�3�f9u���H%   � ���E��a���3�f;�uF�E����u9E�u9E�u	f�E���  f;�uF�E����u9E�u	9E��v����E��}��E�   �E��M���M���~K�M؉M��D��M���	�e� �ʋW��
;�r;�s�E�   �}� �_�tf��m����M��}� ����E��M��}� ����  f��~7�}���x+�E�M��e��������E����?���  �E�f���f��M����  f��yB��������E�t�E��M��}�U��m�������M������H�}�M�u�9E�tf�M�� �  f9E�w�M����� �� � u4�}��u+�e� �}��u�e� ���  f9M�uf�E�F�f�E���E���E��  f;�r#3�3�f9E��E����E�I��   ��� ���M��;f�E�u�f�E��E�E�E��E�f�u��3�f�����e� H%   � ���e� �E��E�U��E��}f�t0����)3�f�� �  f9E�f�B0����$ �B�B �s�����~j_�u������?  3�f�E��E�   �E��]�M��e����؋E������M��]�E�u؅�y2�ށ��   ~(�E�]�M��m�����؋E������N�]�E���؍G�Z�]��E�����   �U��E�u��}ĥ���e��}��e���� ʋU�����֋��4	����U���ȋE���<;�r;�s�F3�;�r��s3�B����tA�Eȍ0�U�;�r;�sAM����ʍ4?�u��u��M������0������C�M��}� �u��E� �K����C���<5}�M��D�;9u	�0K;]�s�E�;]�sCf� �*؀��ˈX�D �E��M�_^3�[��Q���À;0uK;�s��E�;�s�3�f�� �  f9U��@���ʀ��� �P�0�@ ����3���t@��t����t����t����t�� ��   t���˺   #�V�   t#��   t;�t;�u   �   �   �ˁ�   t��   u���^��   t   �3���t��   SVW�   ��t���t   ��t   ��t   �   ��   tǋʾ   #�t;�t;�t;�u `  � @  �    �   _#�^[��   t��   t
;�u �  Ã�@�@�  Ë�U���SVW��}�f�]�3���tjZ��t����t����t���� t����t��   �ˋ��   #ƿ   t$=   t=   t;�u����   ���   #�t��   u��   ���   �é   t��   �}�M����#�#���E;���   ���������E��m���}��]�3���tjZ��t����t����t���� t����t��   �ˋ�#�t(=   t=   t;�u��   ���   ���   ��   t��   u��   ���   ��   t��   �U��3�95T��  ���}��]��E���yj^�   t���   t���   t���   t���   t��   �Ȼ `  #�t*��    t�� @  t;�u��   ���   ���   �@�  #ǃ�@t-�  t��@u��   ���   ���   �E��#E��#��;�u���   ����P�E������Y�]�M�3҄�yjZ��   t����   t����   t����   t���   ��t��   ��#�t$=    t= @  t;�u��   �
��   ��#σ�@t���  t��@u��   ���   ���   ��3ME�� t   �_^[��Q�L$+ȃ����Y��  Q�L$+ȃ����Y��  ��U��QQ�EV�u�E��EWV�E��W  ���Y;�u荖��� 	   �ǋ��J�u�M�Q�u�P���E�;�u����t	P����Y�ϋ����� S�����D0� ��E��U�_^��jhh
��������]܉]��E���u�$����  �	���� 	   �Ë��   ��x;�Rr������  ����� 	   �%����ы����<� S��������L1��t�P��  Y�e� ��D0t�u�u�u�u��������E܉U������� 	   臕���  �]܉]��E������   �E܋U��U�����u�  YË�U���  �F  �`#3ŉE��EV�uW3���4�����8�����0���9}u3��  ;�u�����8������    �<�������  ������S�� S������L8$�����$�����?�����t��u'�M����u贔���  虔���    �ݞ���  �D8 tjj j V������V�>  Y����  ��D���  �i���@l3�9H�� �����P��4����3�;��`  ;�t8�?����P  ����4����� ���3���,���9E�#  ��@�����?������g  ���$���3���
��������ǃx8 t�P4�U�M��`8 j�E�P�K��P�����Y��t:��4���+�M3�@;���  j��D���SP�  �������  C��@����jS��D���P�  ������n  3�PPj�M�Qj��D���QP�� ���C��@�����������=  j ��,���PV�E�P��$���� �4������
  ��@�����0������8���9�,�����  ����� ��   j ��,���Pj�E�P��$���� �E��4�������  ��,�����  ��0�����8����   <t<u!�33Ƀ�
������@�����D��������<t<uR��D����+  Yf;�D����I  ��8�������� t)jXP��D�����  Yf;�D����  ��8�����0����E9�@���������  ����8����T4��D8��  3ɋ�D8���  ��?��� ��D�����   ��4���9M��  ��3�+�4�����H���;Ms&�CA�� �����
u��0���� @F�@F���  rՋ���H���+�j ��(���PV��H���P��$���� �4������C  ��(����8���;��;  ��+�4���;E�l����%  ��?�����   ��4���9M�H  ��@��� ��+�4���j��H���^;MsC��Ή� �����
u�0���j[f��� �����@����@���f�Ɓ�@����  r�����H���+�j ��(���PV��H���P��$���� �4������i  ��(����8���;��a  ��+�4���;E�G����K  ��4�����,���9M�u  ��,�����@��� +�4���j��H���^;Ms;��,�����,���΃�
uj[f���@����@���f�Ɓ�@����  r�3�VVhU  ������Q��H���+��+���P��PVh��  �����;���   j ��(���P��+�P��5����P��$���� �4�����t�(���;�������D���;�\��,���+�4�����8���;E�����?Q��(���Q�u��4����48�����t��(�����D��� ��8��������D�����8��� ul��D��� t-j^9�D���u躎��� 	   ����0�?��D����Ǝ��Y�1��$���� �D@t��4����8u3��$�z����    肎���  ������8���+�0���[�M�_3�^�D����jh�
������]���u�F����  �+���� 	   ����   ��x;�Rr�����  ����� 	   �H����ҋ����<� S�������D0��t�S��  Y�e� ��D0t�u�uS�n������E��認��� 	   貍���  �M���E������   �E�腇��Ë]S�?  YË�U����Bh   �|��Y�M�A��t�I�A   ��I�A�A�A   �A�a �]Ë�U��E���u����� 	   3�]Å�x;�Rr����� 	   �F����ދȃ����� S���D��@]ø@0á�RVj^��u�   �;�}�ƣ�RjP�)|��YY��B��ujV�5�R�|��YY��B��ujX^�3ҹ@0���B��� �����2|�j�^3ҹP0W������ S����������t;�t��u�1�� B���0|�_3�^��
  �=x9 t�m  �5�B�H��YË�U��V�u�@0;�r"���2w��+�����Q豗���N �  Y�
�� V���^]Ë�U��E��}��P脗���E�H �  Y]ËE�� P���]Ë�U��E�@0;�r=�2w�`���+�����P�b���Y]Ã� P���]Ë�U��M�E��}�`�����Q�3���Y]Ã� P���]Ë�U��E��u�����    �W������]Ë@]á`#��3�9�B����Ë�U���SV�u3�W�};�u;�v�E;�t�3��{�E;�t�������v詊��j^�0�������V�u�M���d���E�9X��   f�E��   f;�v6;�t;�vWSV�F�����^���� *   �S���� 8]�t�M��ap�_^[��;�t&;�w �3���j"^�0�x���8]�t��E��`p��y�����E;�t�    8]��<����E��`p��0����MQSWVj�MQS�]�p���;�t9]�j����M;�t�������z�P���;��s���;��k���WSV�E�����[�����U��j �u�u�u�u������]���U��V3�PPPPPPPP�U�I �
�t	���$��u����I ���
�t	���$s���� ^������������U��V3�PPPPPPPP�U�I �
�t	���$��u���
�t���$s�F��� ^�Ë�U����ES3�VW�E�N@  ��X�X9]�E  �]����}襥��э<	���ʋU�e ��ى}����֋u����ϋ��M���U�����։0�x�H;�r;U�s�E   �} �t'�u��e �~;�r��s�E   �} �xtA�H�u�e �7;�r;�s�E   �} �XtA�HM��e� ��ɋ��������މH�M�M�M��X�1�2�u�;�r;�s�E�   �}� �t$�K3�;�r��s3�B�ىH��t
�M�A�M�H�M�M�E�} �X�H�����3�9Xu*�P��E���  ��������������P�;�t܉x�x�� �  u0�H��E���  �����������ʉ�H�x�� �  t�f�M�_^f�H
[��������������Q�L$+����#ȋ�% ���;�r
��Y�� �$�-   � ���U��MS3�VW;�|[;�RsS��������<� S����D0t6�<0�t0�=6u+�tItIuSj��Sj��Sj������3���X���� 	   �`�������_^[]Ë�U��E���u�D����  �)���� 	   ���]Å�x;�Rr� ����  ����� 	   �I����Ջ����� S�����Dt͋]�jh�
����}����������4� S�E�   3�9^u5j
�{���Y�]�9^uh�  �FP�p���u�]��F�E������0   9]�t���������� S�D8P����E��K���3ۋ}j
�=���YË�U��E�ȃ����� S���DP���]Ë�U��Q�=�5�u��  ��5���u���  ��j �M�Qj�MQP����t�f�E�Ë�U���SV�u3�;�t9]t8u�E;�t3�f�3�^[���u�M���^���E�9Xu�E;�t�f�8]�t�E��`p�3�@�ˍE�P�P����YY��t}�E����   ��~%9M| 3�9]��R�uQVj	�p�ذ���E�u�M;��   r 8^t���   8]��f����M��ap��Z��������� *   8]�t�E��`p�����;���3�9]��P�u�E�jVj	�p�ذ���:���뺋�U��j �u�u�u�������]�jh�
�R}��3ۉ]�j�c���Y�]�j_�}�;=�R}T����B9�tE���@�tP��  Y���t�E��|(��B���� P�|���B�4���?��Y��B��G��E������	   �E��}���j����YË�U��SV�u�F�Ȁ�3ۀ�u@�  t9�FW�>+���~,WPV����YP������;�u�F��y����F��N ���_�F�f �^��[]Ë�U��V�u��u	V�5   Y�/V�|���Y��t�����F @  tV�E���P�J  Y��Y��3�^]�jh�
�|��3��}�}�j����Y�}�3��u�;5�R��   ��B��98t^� �@�tVPV�J���YY3�B�U���B���H���t/9UuP�J���Y���t�E��9}u��tP�/���Y���u	E܉}��   F�3��u��B�4�V�S���YY��E������   �}�E�t�E��{���j�~���Y�j����Y���������������̋D$�L$ȋL$u	�D$��� S��؋D$�d$؋D$���[� 3�PPjPjh   @h�������5á�5���t���tP���Ë�U��V�uW�����u�����    �(�����D�F�t8V�����V���N  V����P�~  ����y�����F��tP�2=���f Y�f ��_^]�jh�=z���M��3��u������u�j����    變�������F@t�f �E��Iz���V�?���Y�e� V�<���Y�E��E������   �ԋuV����Y�jh0��y���]���u� ���� 	   ����   ��x;�Rr����� 	   �%����ڋ����<� S�������D��t�S�����Y�e� ��Dt1S�W���YP�����u���E���e� �}� t����M��j��� 	   �M���E������   �E��My��Ë]S����Y�������������U��WVS�M�tM�u�}�A�Z� �I �&
�t'
�t#����:�r:�w�:�r:�w�:�u��u�3�:�t	�����r�ً�[^_�Ë�U��V�uWV����Y���tP� S��u	���   u��u�@Dtj�U���j���L���YY;�tV�@���YP�����u
�����3�V���������� S����Y�D0 ��tW�i~��Y����3�_^]�jhP��w���]���u�1~���  �~��� 	   ����   ��x;�Rr�
~���  ��}��� 	   �3����ҋ����<� S�������D0��t�S�����Y�e� ��D0tS�����Y�E���}��� 	   �M���E������   �E��w��Ë]S�:���YË�U��V�u�F��t�t�v��9���f����3�Y��F�F^]��%��������̋T$�B�J�3��3������30������̋T$�B�J�3��t3���(��0������̋T$�B�J�3��T3�������/������̋T$�B�J�3��43�������/������̋T$�B�J�3��3���0 �/������̋T$�B�J�3���2���� �/������̋T$�B�J�3���2���� �s/������̋T$�B�J�3��2���8�S/������̋T$�B�J�3��2�����3/������̋T$�B�J�3��t2�����/������̋T$�B�J�3��T2���@��.������̋T$�B�J�3��42������.������̋T$�B�J�3��2�����.������̋T$�B�J�3���1���H�.������̋T$�B�J�3���1�����s.������̋T$�B�J�3��1�����S.������̋T$�B�J�3��1���P�3.������̋T$�B�J�3��t1�����.������̋T$�B�J�3��T1��� ��-������̋T$�B�J�3��41���X��-������̋T$�B�J�3��1�����-������̋T$�B�J�3���0����-������̋T$�B�J�3���0���`�s-���T$�B�J�3��0����X-������������h���;��Y����̃=�5 uK��5��t��5�Q<P�B�Ѓ���5    ��5��tV���p���V�jR������5    ^�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           � � � � � � � 
  & B N \ j t � � � � � �   < P X f x � � � � � �  . H V d ~ � � � � � �   ( 2 > P ^ n ~ � � � � � � �           ��        �����7�        Ӟ                            �HR       }   �� �� 0� >�vector<T> too long  --SolidChamfer 2.2, Filip Malmberg 2013--   map/set<T> too long     -DT�!	@      �              �?      @X�0> 04 �0�@�P� �`�����p�����В�����`�p��@�`�p�P��5  �0� �@� �К�    c:\program files\maxon\cinema 4d r12 demo\plugins\solidchamfer2.2\source\sc_modifier.cpp    SolidChamfer Modifier   osolidchamfer   SolidChamferModifier.tif    invalid map/set<T> iterator           �?      �?UUUUUU�?���� � P� �� � � �����c:\program files\maxon\cinema 4d r12 demo\plugins\solidchamfer2.2\source\sc_tool.cpp    ��0> �/00P� @/P/`/p/� �/0� �/�/`0p0�0`� �0�0�0�0 1SolidChamfer    SolidChamfer.tif    Apply Solidchamfer to selected edges.   Apply   Offset  Subdivision     �������������c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_libs\lib_ngon.cpp   $� �p�`9�� �c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_general.h   %s     c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_resource.cpp    #   M_EDITOR        ����MbP?�@��uP� �    c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_baseobject.cpp  ��Бres      �f@��������� �� ���Ш      Y@     @�@��������� �� ���`��@0�@�����P������� ���c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_gui.cpp X�������� �� �����    l�������� �� �����P�`�p����������	 ������Progress Thread 0%  ~   %       c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_file.cpp    c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_basebitmap.cpp      c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_basetime.cpp         �Ngm��C   ����A  4&�k�  4&�kC����Б!�!�    c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_pmain.cpp   �@�c:\program files\maxon\cinema 4d r12 demo\resource\_api\c4d_gv\ge_mtools.cpp    L����� �����(��>�t��>����>���>�Unknown exception   (�l�csm�               �        ��              �?      �?3      3            �      0C       �       ��              fmod         ���d��������p���>�bad exception   K E R N E L 3 2 . D L L     FlsFree FlsSetValue FlsGetValue FlsAlloc    (6�6e+000                 8C      8CX������< 1�
�"�?'���;�< ï&�b�?�,kg��< !J���?ĂeT1��< �1y"�?�z���< �F#�?V���a�< $�
lc�?���x��< �nu���?c�v5��< ����?0��N�< �ߢ�#�?	��"$�< b�md�?�g�Q��< |a7��?�麏��< a��c�?0H_��< �А$�?]U ?�< 8�U�d�?|}}�?�< 5�盧?~+����<  �?)0>�B��< �'HR%�?���I&�< ^:ȅe�?>!ʎ��< sl����?e�cb~q�< �ۧ��?r���ʀ�< F�(&�?Z��n��< '��`f�?4�7j��< ��㚦�?+i��	U�< �oX��?F��.K;�< ��.'�?Yh�ŉ�< 4lkQg�?�;+�U��< 3���?�М	m8�< ��&��?����< �S�(�?Y�=�t< :@�Xh�?,�n@4`�< ��$���?�����< �n��?��9�ܮ�< � �-)�?\�����< �Řwi�?���=�< R�%é�?�f�@��< *�B�?a���w��< G��^*�?�m(�<��< �2;�j�?��P�E�< ����?<�/����< :�T�?Ft����< ͩ+�?N�ibzP�< ��� l�?��  %X�< aY��?]@�_}�< �nL��?����G	�< �1-�?a���(�< U�lm�?iT	�?��< �*̭�?V��*���< w7H-�?��X[F�< �+�.�?X� kn�< E���n�?�T�(�+�< ��U[��?։���< '���?ju!4���< ��-0�?������< Q̙p�?�冿��< �����?���{��< qw�?_W����< �C�1�?'����< I��\r�?��D�c< s�>Ҳ�?������< w*�I�?���n'$�< �2�3�?z���7�< [��>t�?V-Ai��< �����?`�DTb�< �;��?S��.��< TR�*�?)�R���< 2���k�?,�%�ً�< r����?SC?
�< H����?Zxg�f��< �`/-�?����#�< މ7�m�?�w���< 悆a��?_"�C���< lX^��?���@��< �{Х/�?$�8�^�< ]h�Np�?b�X*��< �����?�}�_Ͼ< ��s���?��p�t�< �h�f2�?��$�V�< �4{#s�?U���g
�< ����?��w���< J.����?I�Z��< *�Ow5�?��.@��< ��FHv�?N	����< �!���?�j����< �v(���?��z�"�< i�6�8�? �?!���< <���y�?G��o��< �魺�?�xeF���< �豟��?�G��T��< ��1�<�?V�	ڀ�< ��{�}�?���0���< �����?���a@��< ﶠ��?�0����< ��̯@�?��1�< �3�ā�?��.aU�< !�E���?�I�����< ����?���	���< �j�)E�?O�����< I�W��?W�0�e)�< ��u���?����
T�< �˛��?����?��< �X	J�?!PO79�< �/�Q��?�;�X��< J]���?V:e:���< �Q���?�Wm��`�< b;�SO�?4Td'��< 
Xw���?ЀY��< �L"��?d��ݩS�< _}?��?�T�x�< �[bU�?�\�z#��< ^ɍ��?1����< �N���?�wa���< �����?���N9�< a�X;[�?���Y']�< @ٜ̓�?���E�< VOu��?!S�ÀX�< b- �?C�:���< �|�a�?B�<��$�< �{ɟ��?+X�UG�< m�e��?>Uۊ�< �o]2'�?�� I��< Р�i�?G�����< ��o��? ��Ιn�< 9�[���?�	�|�^�< ����.�?�>oj��< .�_�p�?1S���< �X����?����l�< �~���?o.x���< %3d�?����{ = 4 ��L�?�V!�= b�#��?��@g	= a��?G��z	= �]ư�?���6�= o�JV�?J�� �b= '4��?/��t�>�< w���?a�`����< �_��?a�	�e= ��F``�?/�f	= #&��?�5SmT4�< W�� ��?R�z��<  ъ�(�?���vY�< ���k�?p�Y�.= �y���?�8�'���< Ku�C��?j��<{= 2�<�5�?��ýd	= ��x�?�"a��= @�ic��?�%�[�9= �����?kR�F��< �6D�C�?ş
ܬ_�< 5��Z��?ȡ�k*= ���3��?�*+xi(�< �G�&�?��r
ly= :��3S�?z
�j�< �[��?��'����< ;!���?h����= �<��?���:��< ��sd�?��3�= �?	��?{�!m�B�< <>����?�*�2 = ����2�?cM�yoG= V��sw�?8K��$�< ��}��?C�l���< Ϲ���?�-��< '���F�?ɕ���{�< �$�R��?܊�)B��< �#���?������< ��c�?? ��~��< ���F]�?���&��= �		/��?94��E�< ?T9��?9*��)�< l?�e/�?�B6�!F= u0w�u�?�M�떐= �k`(��?������< 4�=��?Kp��= G"�zI�?$�}Tw5�< �[��?ߪ��b�< �Ka��?aF7�= Vj��?�T��y�< R߂�e�?M]-��e�< $�[��?3����< Ễ���?��QZo�= n��<�?1-
I�x�< f�	���?I��]�= ��O���?���x�= �#$�?�nz��= �) �]�?����h��< �'�7��?y]h�= �Yg��?�S�c�< b}��?��$ګ= ;�ђ@�?OD���)= ���=e�?:Q�]D\�< ��� ��?FnH�AY�< "�ۮ�?�)Bp�= )R�Q��?��{���< �L��0�?�U��< d�N{�?���c�1= f��k��?iO��)= ��m��?�
��R = l[��]�?�$Ŝi= w/�d��?���C�= �(�O��?u��1��= ��/�D�? �&= �� ���?i�C1]�< Ei��?X�=g��< P�~0�?Y;���=  ]��?���m��< �����?�A�8�y�< �7�l �?S6���= =.�q�?+`���= �����?���%!5= �o�h�?�y���= i�Q�i�?v�7���= �Խ�?dDR޸;= nl���?b*t#�= x�A@h�?�����= ZmI���?�oP�@= ��Y��?��Ͽ	= �n�?u�И?�= %�k��?ZEM-'^= DT!�?:Z��n== ��0|�?�O���= ���*��?m}I�{= �eP5�?+�}ZI= �Q����?�^oc;�< '��?
u�/r��< ���S�?�i���1= �q���?/����= {�ss�?VV&�= �#�k~�?[��	�< �����?vB���< 6��#M�?��!��< 
��?q_�w#�< ����"�?ұ��R��< �����?k=�C= �B� �?��_���< u���r�?�y���= Dw�b��?�(,xn�< <"Q/�?���q�q)= �o\l�?�)���T&=  7a��?��L�< �?|6��?�������?#�DZ9��?������?��/�.��?>6)}���?, �,��?��؏��?M�����?��x%q��?�� ����?/x�bJ��?Ȉb����?�uÏ��?(Z����?��t����?{}�2F��?�������?_�2��?>�T�^��?�u	���?�����?4t��d��?��Z���?(�	��?WI�Y��?�d���?�{�����?|��:��?�S9���?���s���?���
��?����K��??�����?l�.���?�Z�3��?��;E<��?�fSOs��?�J�Q���?�z�L���?�@��?{yK+;��?ãjh��?��F���?-(�����?�n�����?@��F��?����)��?�P�J��?C��Si��?�^����?�B����?i|e���?�������?�� ���?�a�k���?c����?X�!��?89�l!��?fh�+��?��3��?)Ao
:��?�1(>��?2:@��?>�?@@��?"I�r���?6��4���?�@Û��?����?765@Z��?�&+-��?w�'����?��Q���?�Gp�t��?�2�&��?X��9Ш�?B�q��?/�?�
��?v�ɛ��?��Mj$��?�3����?�s����?b里��?V�����?%S��?V��ѩ��?ߖ%@���?�U>��?2�,|��?�ܜm���?V��kށ�?9�?�I�@|�?��P3y�?�?}>v�?��H|As�?#�<p�?_0.m�?t���j�?���f�?�����c�?�3)�`�?��i]�?�� F)Z�?�2V�V�?��f\�S�?B?}4P�?���V�L�?{�fI�?uS�E�?|�ǩuB�?1�<��>�?�(��b;�?�탿�7�?�]o�-4�?P�h�0�?�H�,�?�:5�)�?Iٓ\%�?f,��!�?갸%��?N���?$�k��?�oay�?*���?��?Y
�?���$�?�?�(�?���a���?�9y����?99R��?%��R���?F�����?��@�I��?j �T��?�0<��?2j���?�p�~���?,�L��?@�_�o��?7�����?�'�����?�VG��?�D<xZu�?`\@��j�?)]G�q`�?L�c�U�?�Jup�J�?CY���?�?� X7�4�?�T��)�?KB	�0�?&D��?lU����?�E0d��?KYC ��?�:����?@М����?��L���?#�e�m��?-Fգ��?�DT����?�W�㗖�?*�MU��?�z��{�?�l�Un�?
Q-��`�?>�ұR�?V�D��D�?oW�sg6�?U��J(�?>��t�?2̄λ
�?�1_����?$*2���?[��ێ��?N��)��?���V���?l$G~ٮ�?��+6��?�tF4؎�?��,�~�?����"n�?<�փ]�?|ߠ�L�?l6���;�?6*��*�?�|�59�?��:��?H�K����?s7��?��I-���?�$z����?�9\���?��>|.~�?�-��W�?�^\sY0�?:Rp�7�?m�bzA��?G�4's��?I�y�Ȋ�?%��=_�?�C\�2�?�O��u�?�m��.��?�M����?���n�w�?KK�'�F�?��l^�?:��" ��?��Ѭ�?��}6lw�?�:�@�? 7Z8>	�?$�� f��?e')lW��?zD@	[�?���jq�?�P J���?F���<��?�Q'J�`�?x��e_�?* Aӱ��?�"�Sr��?xw��N�?k��$��?
�S/���?��yx|o�?P�6 d!�?ZyrI��?�����?��Ӳ�*�?
T�����?���!�z�?��{��?��0�V��?�8I�^�?��A;��?���wC��?�JG7�&�?�'un�?���)��?m���y��?������?��|�ȕ�?,"��Q��?�/��b�?PV3� 2�?�S����?p����?V�a��"�?�Tl��?Pq�j��?��Y��?p�,�?�l"։�?cY�����?\3&��<-DT�!�?\3&���-DT�!	�\3&��<-DT�!	@       �           �����   �����    ���                UUUUUUſ333333���m۶mۦ�颋.��?333333�?�q�q�?UUUUUU�?O��N�đ?�m۶mۦ?$rxxx��?�������?�������     ���      �?      �?       �9��B.�@  ׽2b      �              �7       ���5�h!����?      �?            �?5�h!���>@�������             ��      �@      �        CorExitProcess  m s c o r e e . d l l         �         �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       �  �       � �       � �          	   �      r u n t i m e   e r r o r        
     T L O S S   e r r o r  
   S I N G   e r r o r  
     D O M A I N   e r r o r  
     R 6 0 3 3  
 -   A t t e m p t   t o   u s e   M S I L   c o d e   f r o m   t h i s   a s s e m b l y   d u r i n g   n a t i v e   c o d e   i n i t i a l i z a t i o n 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .   I t   i s   m o s t   l i k e l y   t h e   r e s u l t   o f   c a l l i n g   a n   M S I L - c o m p i l e d   ( / c l r )   f u n c t i o n   f r o m   a   n a t i v e   c o n s t r u c t o r   o r   f r o m   D l l M a i n .  
     R 6 0 3 2  
 -   n o t   e n o u g h   s p a c e   f o r   l o c a l e   i n f o r m a t i o n  
     R 6 0 3 1  
 -   A t t e m p t   t o   i n i t i a l i z e   t h e   C R T   m o r e   t h a n   o n c e . 
 T h i s   i n d i c a t e s   a   b u g   i n   y o u r   a p p l i c a t i o n .  
     R 6 0 3 0  
 -   C R T   n o t   i n i t i a l i z e d  
     R 6 0 2 8  
 -   u n a b l e   t o   i n i t i a l i z e   h e a p  
         R 6 0 2 7  
 -   n o t   e n o u g h   s p a c e   f o r   l o w i o   i n i t i a l i z a t i o n  
         R 6 0 2 6  
 -   n o t   e n o u g h   s p a c e   f o r   s t d i o   i n i t i a l i z a t i o n  
         R 6 0 2 5  
 -   p u r e   v i r t u a l   f u n c t i o n   c a l l  
       R 6 0 2 4  
 -   n o t   e n o u g h   s p a c e   f o r   _ o n e x i t / a t e x i t   t a b l e  
         R 6 0 1 9  
 -   u n a b l e   t o   o p e n   c o n s o l e   d e v i c e  
         R 6 0 1 8  
 -   u n e x p e c t e d   h e a p   e r r o r  
         R 6 0 1 7  
 -   u n e x p e c t e d   m u l t i t h r e a d   l o c k   e r r o r  
         R 6 0 1 6  
 -   n o t   e n o u g h   s p a c e   f o r   t h r e a d   d a t a  
   R 6 0 1 0  
 -   a b o r t ( )   h a s   b e e n   c a l l e d  
     R 6 0 0 9  
 -   n o t   e n o u g h   s p a c e   f o r   e n v i r o n m e n t  
   R 6 0 0 8  
 -   n o t   e n o u g h   s p a c e   f o r   a r g u m e n t s  
       R 6 0 0 2  
 -   f l o a t i n g   p o i n t   s u p p o r t   n o t   l o a d e d  
            ��   X�	    �
   ��   `�    �   ��   `�   ��   ��   0�   ��   p�   0�   h�     �!   �x   ��y   ��z   ���   ���   ��M i c r o s o f t   V i s u a l   C + +   R u n t i m e   L i b r a r y     
 
     . . .   < p r o g r a m   n a m e   u n k n o w n >     R u n t i m e   E r r o r ! 
 
 P r o g r a m :           �      ��      �                       �  �  ��  �  ��       ���Iq��I�`B�`B��Y���n�Y���n��tan cos sin modf    floor   ceil    atan    exp10   acos    asin    log log10   exp pow �������             ��      �@      �         Complete Object Locator'    Class Hierarchy Descriptor'     Base Class Array'   Base Class Descriptor at (  Type Descriptor'   `local static thread guard' `managed vector copy constructor iterator'  `vector vbase copy constructor iterator'    `vector copy constructor iterator'  `dynamic atexit destructor for '    `dynamic initializer for '  `eh vector vbase copy constructor iterator' `eh vector copy constructor iterator'   `managed vector destructor iterator'    `managed vector constructor iterator'   `placement delete[] closure'    `placement delete closure'  `omni callsig'   delete[]    new[]  `local vftable constructor closure' `local vftable' `RTTI   `EH `udt returning' `copy constructor closure'  `eh vector vbase constructor iterator'  `eh vector destructor iterator' `eh vector constructor iterator'    `virtual displacement map'  `vector vbase constructor iterator' `vector destructor iterator'    `vector constructor iterator'   `scalar deleting destructor'    `default constructor closure'   `vector deleting destructor'    `vbase destructor'  `string'    `local static guard'    `typeof'    `vcall' `vbtable'   `vftable'   ^=  |=  &=  <<= >>= %=  /=  -=  +=  *=  ||  &&  |   ^   ()  ,   >=  >   <=  <   /   ->* &   +   -   --  ++  *   ->  operator    []  !=  ==  !   <<  >>  =    delete  new    __unaligned __restrict  __ptr64 __eabi  __clrcall   __fastcall  __thiscall  __stdcall   __pascal    __cdecl __based(         �����������������������������|�x�t�p�l�h�\�X�T�P�L�H�D�@�<�8���4�0�,�(�$� ���������� ���������������������������d�D�$����������`�8���� �������������l�D����������d�8��������������p�H H : m m : s s     d d d d ,   M M M M   d d ,   y y y y   M M / d d / y y     P M     A M     D e c e m b e r     N o v e m b e r     O c t o b e r   S e p t e m b e r   A u g u s t     J u l y     J u n e     A p r i l   M a r c h   F e b r u a r y     J a n u a r y   D e c   N o v   O c t   S e p   A u g   J u l   J u n   M a y   A p r   M a r   F e b   J a n   S a t u r d a y     F r i d a y     T h u r s d a y     W e d n e s d a y   T u e s d a y   M o n d a y     S u n d a y     S a t   F r i   T h u   W e d   T u e   M o n   S u n   HH:mm:ss    dddd, MMMM dd, yyyy MM/dd/yy    PM  AM  December    November    October September   August  July    June    April   March   February    January Dec Nov Oct Sep Aug Jul Jun May Apr Mar Feb Jan Saturday    Friday  Thursday    Wednesday   Tuesday Monday  Sunday  Sat Fri Thu Wed Tue Mon Sun GetProcessWindowStation GetUserObjectInformationW   GetLastActivePopup  GetActiveWindow MessageBoxW U S E R 3 2 . D L L     ( n u l l )     (null)         EEE50 P    ( 8PX 700WP        `h````  xpxxxx          _nextafter  _logb   _yn _y1 _y0 frexp   fmod    _hypot  _cabs   ldexp   fabs    sqrt    atan2   tanh    cosh    sinh                                                                                                                                                                                                                                                                                          ( ( ( ( (                                     H                � � � � � � � � � �        � � � � � �                           � � � � � �                                                                                                                                                                                                                                                                                                               h ( ( ( (                                     H                � � � � � � � � � �        ������      ������                                                                      H                                      �������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@abcdefghijklmnopqrstuvwxyz[\]^_`abcdefghijklmnopqrstuvwxyz{|}~���������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������� 	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`ABCDEFGHIJKLMNOPQRSTUVWXYZ{|}~��������������������������������������������������������������������������������������������������������������������������������	
 !"#$%&'()*+,-./0123456789:;<=>?@ABCDEFGHIJKLMNOPQRSTUVWXYZ[\]^_`abcdefghijklmnopqrstuvwxyz{|}~ 1#QNAN  1#INF   1#IND   1#SNAN  C O N O U T $   ������  �����EEE���  00�P��  ('8PW�  700PP�    (����   `h`hhhxppwpp           H                                                           `#��   RSDSp���(K�E�<y�   C:\Program Files\MAXON\CINEMA 4D R12 Demo\plugins\SolidChamfer2.2\obj\SolidChamfer_Win32_Release.pdb                  D�           T�`�|�             ����    @   D�         ����    @   ��           ��|�               ������    8        ����    @   ��P         ����    @   �           ���               ,�<�����    h        ����    @   �            � l�           |���<�����    �        ����    @   l�            � ��           ������4�    �        ����    @   ���        ����    @   �           (���4�    �         ����    @   P�           `�4�               x�����    �        ����    @   h�            !��           ��������    !       ����    @   ��            ��    ,!        ����    @   ��            L!8�           H�T��    L!       ����    @   8�            t!��           �����    t!       ����    @   ��            �!��           �����    �!       ����    @   ��            �!�           ,�4�    �!        ����    @   �            �!d�           t����    �!       ����    @   d�            P �            � P�            �!��           ����4�    �!       ����    @   ��            "$�           4�<�    "        ����    @   $�            � �            ,"��           ������4�    ,"       ����    @   ��            H"��           ����    H"        ����    @   ��            `"�           (�0�    `"        ����    @   �            |"`�           p�x�    |"        ����    @   `�            �"��           �����    �"       ����    @   ��            �"��           ��    �"        ����    @   ��            �"<�           L�X�|�    �"       ����    @   <�            �"��           ����X�|�    �"       ����    @   ��            #��           ����X�|�    #       ����    @   ��             ��            <#<�           L�T�    <#        ����    @   <�            �#��           ����|�    �#       ����    @   ��    4� >�   �, �7 �� Т � � 0� P� p� �� �� У � � 0� P� p� �� �� Ф � � 0� P� p� ��                               X�   d���          ����       @          ����       7�            � ����    ����                  ��"�   ��   ��                            �' ����    ����                  ��"�   �   �                            y( ����    ����                  L�"�   \�   l�                            �) ����    ����                  ��"�   ��   ��                            �* ����    ����                  ��"�                                    �0 ����    ����                  T "�   d    t                             �_ ����    ����                  � "�   �    �                             �` ����    ����                  "�      $                            n ����    ����                  \"�   l   |                            t ����    ����                  �"�   �   �                            {� ����    ����                  "�      ,                            K� ����    ����                  d"�   t   �                            � ����    ����                  �"�   �   �                            u� ����    ����                  "�   $   4                            5� ����    ����                  l"�   |   �                            ݝ ����    ����                  �"�   �   �                            �� ����    ����                  "�   ,   <                            �� ����    ����                  t"�   �   �                            Y� ����    ����                  �"�   �   �                            e� ����    ����                  $"�   4   D                            �� ����    ����                  |"�   �   �                            �� ����    ����                  �"�   �   �                            �� ����    ����                  ,"�   <   L                    �"    ����       f�    a�    �   ����    �"    ����       ��    a�    �   ����    #    ����        �����    ����    ����    ��    ����    ����    ����!�2�    ����    ����    ����    h�    ����    ����    ����    ��    ����    ����    ����    7�    �������    ����    ��������@           ������    ����                  �"�   �   �                   ����    ����    ����    ��    i�r�����    ����    ��������    ����    ����    ����y�}�    ��    �   ���    �#    ����       p�    ����    ����    ����    ������    ������    ����    ����    T�����    `�����    ����    ����u�y�    ����    ����    ��������    ����    ����    ����    i    ����    ����    ����    �+    ����    ����    ����    �0    ����    ����    ����    ~3    ����    ����    ����    P7    ����    ����    ����    �C    ����    ����    ����;ENE    ����    ����    ����3`O`    ����    ����    ����    ��    ����    ����    ����    a�    ����    ����    ����    ��    ����    ����    ����    ՜    ����    ����    ����    _�        +�����    ����    ����    ��    ����    ����    ����    ��    ����    ����    ����    f��         *  �                     � � � � � � � 
  & B N \ j t � � � � � �   < P X f x � � � � � �  . H V d ~ � � � � � �   ( 2 > P ^ n ~ � � � � � � �       �RaiseException  RtlUnwind �GetCurrentThreadId  � DecodePointer �GetCommandLineA �HeapAlloc GetLastError  �HeapFree  � EncodePointer IsProcessorFeaturePresent �TlsAlloc  �TlsGetValue �TlsSetValue �TlsFree �InterlockedIncrement  GetModuleHandleW  sSetLastError  �InterlockedDecrement  EGetProcAddress  �TerminateProcess  �GetCurrentProcess �UnhandledExceptionFilter  �SetUnhandledExceptionFilter  IsDebuggerPresent �Sleep ExitProcess oSetHandleCount  dGetStdHandle  �InitializeCriticalSectionAndSpinCount �GetFileType cGetStartupInfoW � DeleteCriticalSection GetModuleFileNameA  aFreeEnvironmentStringsW WideCharToMultiByte �GetEnvironmentStringsW  �HeapCreate  �HeapDestroy �QueryPerformanceCounter �GetTickCount  �GetCurrentProcessId yGetSystemTimeAsFileTime %WriteFile GetModuleFileNameW  �HeapSize  9LeaveCriticalSection  � EnterCriticalSection  rGetCPInfo hGetACP  7GetOEMCP  
IsValidCodePage �HeapReAlloc ?LoadLibraryW  -LCMapStringW  gMultiByteToWideChar iGetStringTypeW  fSetFilePointer  �GetConsoleCP  �GetConsoleMode  �SetStdHandle  $WriteConsoleW � CreateFileW R CloseHandle WFlushFileBuffers  KERNEL32.dll              �HR    r          h l p 0� �   SolidChamfer.cdl c4d_main                                                                                                                     �    .?AVbad_alloc@std@@ �    .?AVexception@std@@ �    .?AVNodeData@@  �    .?AVBaseData@@  �    .?AVObjectData@@    �    .?AVSC_Modifier@@   �    .?AVSC_ToolDialog@@ �    .?AVSubDialog@@ �    .?AVGeDialog@@  �    .?AVToolData@@  �    .?AVSC_Tool@@             @   �    .?AVGeSortAndSearch@@   �    .?AVTranslationMapNewSearch@@   �    .?AVTranslationMapSearchN@@ �    .?AVTranslationMapSearch@@  �    .?AVNeighbor@@  �    .?AVDisjointNgonMesh@@  �    .?AVGeModalDialog@@ �    .?AVGeUserArea@@    �    .?AViCustomGui@@    �    .?AVC4DThread@@ �    .?AVGeToolNode2D@@  �    .?AVGeToolDynArray@@    �    .?AVGeToolDynArraySort@@    �    .?AVGeToolList2D@@  �    .?AVlogic_error@std@@   �    .?AVlength_error@std@@  �    .?AVout_of_range@std@@  �    .?AVtype_info@@             N�@���Du�  s�  acos            sqrt            �    .?AVbad_exception@std@@ ��������        /?/?/?/?/?/?/?/?/?/?        �����
                                                                                           	               	      
                                                !      5      A      C      P      R      S      W      Y      l      m       p      r   	         �   
   �   
   �   	   �      �      �   )   �      �      �      �      �      �      �                    ?                                                                                                                                                                                                                                                                                            C       ������������������������������|�x�t�p�l�h�d�`�\�X�T�L�@�8�0�p�(� ������������������	         ��������������p�`�P�<�(�������������������������������t�h���\�P�@�,���������������                                                                                           �&            �&            �&            �&            �&                              �/        P���X��&@(                                                                                                                                                                                                                                                                                                                                        abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                                                                                                                                                                                                                                                                                                                                       abcdefghijklmnopqrstuvwxyz      ABCDEFGHIJKLMNOPQRSTUVWXYZ                                                                                                                                      )�  `�y�!       ��      ��      ����    @~��    �  ��ڣ                        ��      @�      �  ��ڣ                        ��      A�      �  Ϣ� ��[                 ��      @~��    Q  Q�^�  _�j�2                 ������  1~��     �            ����            p�`��&         8�   <�   ,�   0�   D�   <�!   4�   $�   �   �   ,�   $�   ��   ��    ��   �   ��   �   ��   �   �   �   ��   ��"   ��#   ��$   ��%   ��&   ��      �      ���������              �       �D        � 0         .   .   �/�B�B�B�B�B�B�B�B�B�/�B�B�B�B�B�B�B�/P�R�T�   ���5      @   �  �   ����                     �B    �B                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                .                   �@         �@         �@        @�@        P�@        $�@       ���@        ��@     ���4@   ������N@ �p+��ŝi@�]�%��O�@q�וC�)��@���D�����@�<զ��Ix��@o�����G���A��kU'9��p�|B�ݎ�����~�QC��v���)/��&D(�������D������Jz��Ee�Ǒ����Feu��uv�HMXB䧓9;5���SM��]=�];���Z�]�� �T��7a���Z��%]���g����'���]݀nLɛ� �R`�%u    �����������?q=
ףp=
ף�?Zd;�O��n��?��,e�X���?�#�GG�ŧ�?@��il��7��?3=�Bz�Ք���?����a�w̫�?/L[�Mľ����?��S;uD����?�g��9E��ϔ?$#�⼺;1a�z?aUY�~�S|�_?��/�����D?$?��9�'��*?}���d|F��U>c{�#Tw����=��:zc%C1��<!��8�G�� ��;܈X��ㆦ;ƄEB��u7�.:3q�#�2�I�Z9����Wڥ����2�h��R�DY�,%I�-64OS��k%�Y����}�����ZW�<�P�"NKeb�����}�-ޟ���ݦ�
    ����                                                                                                               (   00Q0�0�0�5�5�566N6�96=H=�=�=    D   �1�1�12F2�2�2>3V3�3�3T5	6�6�6�6�6v7�788�89)9�9�9:�:N;> 0  �   60H0�0�0�1�1$2Q2t2�2�2�3�3444G4M4h44�4�4�4�4�455#555U5w5�5�5�56[6t6�6�67#7<7k7�7#8�9�9:;:�:�:8;C;L;P;T;X;b>i>�>�> @      1V3:!:::E:^:i:�:�:j;�> P     z6�8�:
=&?8?�?�?�?   `     0(0�0&3v5.=v=�= p     �3�3B4G4�7�8�=   �     �0�5 �  L   }3�3�3�3�3�344�67�7�7�7�7r8w8�8�8B9G9�9�9�:�:V=h=>>&>8>�>�>)?   �  x   �1&585�5�59!9e9l9�9�9�9�9�9�9	::#:5:>:P:b:�:�:�:�:;4;l;�;<=<�<�=�=>.>@>R>d>�>�>�>�>�>?!?3?S?z?�?�?�?�?�?�? �  L   0W0�0�0�0�0�0141Y1~1�1�1�1E2c22�2�2�3�4�6�627R8_9j9�9:;�=�=F?]?   �     0p9 �     H1P:c??�?�?�?�?�?   �  @   0/0�0�0�0�0�1�1f2�4�4�5�5&888Y89(9�9�9:I;V=h=>>6>   �  \   5!5?5a5�5�5�5�5c6u6�6�6Y7u7�7�7Y8|8�8�8�8�8959�9�9L:q:�:�:_;t;�;�;�;�;</<T<t<�<�<   @   �9�9�9%:e:�:�:5;u;�;�;<U<�<�<=E=�=�=�=">R>�>�>�>5?�?�?  l   0U0�0�0%1�1�1�3�3�4�6X7\7`7d7h7K8Y8x8�89&9K9S9: :Q:_:�:�:�;�;�;<p<~<�<�<�=�=�=>E>�>�>?E?�?�?     p   0U0�0�051�1�1%2u2�23e3�34U4�4�455�5�5%6u6�67e7�78U8�8�8E9�9�95:u:�:;E;�;�;5<�<�<%=u=�=%>u>�>?�?   0 �   0U0�0�0E1�1�152�2�2%3u3�3%4e4�45U5�5�5Q6�6�6A7�7�7A8�8�8A9�9�9�9�9�9:4:d:�:�:�:�:$;D;t;�;�;�;$<D<d<�<�<�<�<==1=D=a=q=�=�=�=�=>A>Q>d>�>�>�>?$?A?Q?a?t?�?�?�?�? @ �   040_0�0�0�0�01141T11�1�1�1$2J2t2�2�2�2�2343T3t3�3�3�34W4�4�45T5�5�5�56A6a6t6�6�6�6�67$7D7d7�7�7�7�7&8D8a8�8�8�8�8949T9�9�9�9�9:":6:F:t:�:�:�:�:;@;T;d;�;�;�;�;<M<[<n<�<�<�<�<�<==2=B=d=�=�=�=�=>>D>\>�>�>�>�>�>	??&?T?l?�?�?�?�?   P L   00'060d0�0�0�0�0�01D1m1�1�1�1�1�1$2D2d2�2�2�2�2343T3q3�3�3�3�3444T4t4�4�4�4�4545T5q5�5�5�5�5�56!6D6Y6k6t6�6�6�6�6�6�67a7h7�7�78:8I8t8}8�8�8�8�8�8�8�899(9F9e9w9�9�9�9�9�9:":/:G:Y:k:}:�:�:�:�:�:;;4;F;X;a;;�;�;�;�;�;$<2<?<W<i<{<�<�<�<�<�<�<=(=D=V=h=q=�=�=�=�=�=>>->N>d>�>�>�>�>�>�>�>	??-???H?f?�?�?�?�?�?�?   ` �   00/0P0f0�0�0�0�0�0�01 121D1M1k1�1�1�1�1�12!2A2�2�2�2�2�2�2303A3J3]3�3�3�344,4>4d4�4�4�455$5}5�5�5�5�5�5626O6�6�647I7k7�7848T8t8�8�8�8919T9�9�9�9�9$:T:�:�:�:2;Q;q;�;�;�;<1<Q<q<�<�<�<=4=d=�=�=�=�=>4>a>�>�>�>�>??4?�?�? p �   !040T0�0�0�01!1Q1t1�1�1�12$2q2�2�2�23D3d3�3�34[4�4�4�4�45D5q5�5�5�5�5�5*6D6�6�6�6
7T7t7�7P8�8�899=9q9�9�9�9:?:�:�:�:�:(;Y;�;$<4<a<�<�<�<='=E=d=�=�=�=�=$>D>t>�>�>�>�>A?d?�?�?�? � �   0$0D0�0�0�01Q1t1�1�1�12>2Z2v2�2�23#3Q3q3�3�3�3�3464X4n4�4�4�4�45(5g5�5�5�5�56+6@6\67.7z7�7�7�7�7D8W:�<=d=w=�=�=�=4>O>   � �   0000K0P0�0�0�0�0�01$1D1a1t1�1�1�1*3<3N3�3P4W4^4e4l4s4z4�4�4�4�4�4�4�4�4�4�4�5�5616T6t6�6�6�6�67D7d7�7�7�7�78;8a8�8"9�9�9�9:2:�:�:-;�;�;G<�=�=�=�=�=�=�=�=^>j>v>�>�>Q?q?�?�? � �   0T0�0�01$1D1d1�1�1�1�12$2T2t2�2�2�23D3d3�3�3�34?4a4�4�4�45A5a5�5�5�5�56!6A6a6�6�6�6�67!7A7a7�7<8h8�8�8�89W9%:*:5:X:b:�:�:�:�:!;T;�;�;<D<k<�<�<
=6=K=t=�=�=+>k>�>�> ?d?�?�?�?�? � �   0'0V0m0�0�0�0121Q1p1�1�1�1222Q2�2�2�2�23'3g3�3�3�3�3*4�4�4%5~5�56[6�6�6�6;7|7�7�7�7<8V8�8�89!9x9�9�9�94:�:;U;_;�;�;<-<Q<c<v<�<�<�<-=~=�=>Q>�>�>�>"?[?w?�?�?�?�? � x   !0Z0z0�0d1�1�1P2�2�203�3�3C4�4�4C5�56c6�6#7�7�7C8�8 9S9�9:y:�:;�;�;0<`<�<�<�< =P=�=�=�==>a>�>�>�>?>?z?�?�?   � �   K0�0�0.1n1�1�1242q2�2�23T3�3�34%4>4d4�455:5E5[5x5�5�5�5H6d6�67�7&8x8|8�8�8�8�8�8�8�8�8{9�9�9�9�9�9�9�9�9�9�:�:�:�:;";>;a;�;�;�;�;<4<d<�<�<�<=D=�=�=�=>1>Q>k>�>�>$?D?d?�?�?�? � �   0D0t0�0�0�0�0�01#171T1d1�1�1�1�1�1�12"2?2K2V2t2�2�2!3A3d3�3�3 4p4�4�4�4F5t5�5�56T6n67D7�7�7�7�7`8�8�8�8�8�9�9X:�:�:�:�:�:�:�:A;�;�;�;�;
<<D<d<�<(=�=	>4>d>�>�>�>?5?O?l?   � �   0C0a0�0�0�01&1:1O1t1�1�1!2X2]2i2�2�2�2�2$3!4_4�4�4�4�4�45@5a5}5�5�5�5
6.6G6`6�6�6�6 7'7q77�7�7�7�7�78,8J8e8�8�8�8 9V9�9�9~:�:�:�:#;M;t;�;�;<4<�<�<�<�<�<�<='=G=[={=�=�=�=�=�=�=>/>A>T>e>x>�>�>�>   �   p0x0�0�1�12d2�293�34q4�4�4595e5�5�5�6�6t7�7�7�7�7�7�78 828F8c8�8�8�8	9)9=9Y9�9�9�9�9::2:E:Y:k:}:�:�:�:�:�:;);@;v;�;�;�;�;L=S=�=�=�=>1>Q>d>�>�>�>�>$???_?r?�?�?�?�?    �   $0d0�0�0�0�0141T1�1�1�1�1!2D2�2�2�2�23$3D3d3�3�3�3�34444T4t4�4�4535�5�516W6�6(7J7m7�7
8-8�8�8�8N9n9�9:,:T:�:�:�:�;�;�;c<�<�<3=\=�=�=>3>�>?G?�?�?   �   !0G0�0�0!1�12,2T2�2�23~3�3�34a4�4<5d5�5�5�5�5�56+6P6t6�6�67!7D7d7�7�7�7�7!8R8p8�8�8�8�89W9f9�9�9�9:!:D:�:�:�:�:;1;T;�;�;�;�;�;$<T<�<�<�<�<�<=%=g=�=�=�=7>r>�>�>?t? 0 �   040141T1�1�1�12D2t2�2�2�2$3�3�3444"4)40474>4H4R4Y4`4g4n4u4|4�4�4�4�4�4�4�45=5N5_56�6�7�7�7�7848T8�8�8�8�89&9T9t9�9 @    �0�0�0�0�0�01141E1S1q1�1�1�1�12242L2`2p2�2�2�2�2�2�2343L3`3o33�3�3�3�3�344A4Q4d4�4�4�4�45&545G5d5�5�5�56!646T6�6�6�6�6�6747T7t7�7�7�7�7�78$8D8d8�8�8�8�89959d9~9�9�9�9�9:-:D:�:�:�:�:�:;g;�;�;�;�;�;�;H<�<�<�<�<=D=d=�=�=�=�=>$>D>a>t>�>�>�>�>?1?D?_?m?{?�?�?�?�?�?   P (   0!0D0d0�0�0�0�0�0�0�01/1=1K1Z1l1�1�1�1�1242T2t2�2�2�2 33-3W3i3�3�3�3�3�3444T4t4�4�4�4�4�4�4545N5b5q5�5�5�5�5�56,6=6K6b6w6�6�6�6�6�677&7q7�7�7�7�7�78$8D8d8�8�8�8�89$9D9d9�9�9�9�9:$:D:d:�:�:�:�:;@;d;�;�;�;�;<$<D<d<�<�<�<�<=$=D=d=�=�=�=�=>$>D>d>�>�>�>�>�>?1?D?a?q?�?�?�?�?�? ` �   
00D0d0�0�0�01"1�1�1�1T2t2�2�2�2�2�243Q3d3w3�3�3�4�4�4%5e5�5�5%6u6�6�6�657�7�78U8�8�8959�9�9:E:�:�:;5;u;�;�;<e<�<�<5=u=�=�= >>$>E>�>�>?R?�?�?   p �   %0r0�0�0191C1p1u1�1�1�1292u2�2�2�2U3y3�3�3464_4�4�45(5G5h5�5�56T6q6�6�6�67D7q7�7�7�7�7848d8�8�8�8�8949a9t9�9�9�9:4:d:�:�:�:�:4;t;�;�;�;�;<4<T<�<�<�<�<q=�=�=�=>$>�?   � �   
00@01&1�2�2�2$3T3t3�3�3�3�3�3444d4�4�4�4�4�4!5D5a5�5�5�5�56�6,7�7�7�799&9�9�9�9B:�:�:(;6;g;�;�;W<�<�<�<�<�<8=X=v=�=�=�=u>�>�>�>�>�>�>�>?<?a?t?�?�?�?�?   � �   "0>0H0S0X0�0�0�0�0)1Q1q1�1�1�1U2r2�2�2�2�23$3D3a3q3�3�3�3�3�3�3444T4t4�4�4�4�45D5d5�5�5�5�56$6D6�6�6�6�6�67!7?7a77�7�7�7818T8t8�8�8�8�89$9A9T9t9�9�9�9:B:u:�:E;�;�;<U<�<�<2=b=�=�=5>u>�>�>R?�?�?   � |   20b0�0�0121e1�1282L2\2z2�2�2%3u3�34U4�4�4E5�5�5"6b6�6�627x7�728x8�829u9�9:e:�:;R;�;<�<=U=�=�=>e>�>?E?�?�?   � �   50�0�01e1�12e2�2�23-3e3�3�354�4�4%5u5�5%6�6�67U7�7�7%8e8�89^9�9�9:]:�:�:,;;�;<\<�<==D=Q=W=�=�=�=�=�=>>4>8><>@>D>H>Q>t>�>?D?�?�? � t   h0y0�3M4]4�5�5U6�6�6�6�6�6�6M7�78$8�8�8�9F:�:�:�: ;+;:<x<�<�<�<�<�<=F=�=>>H>a>�>�>:?l?�?�?�?�?�?�?�?�?   � 0  0000 0$0(0,000z0�0�0�0�0�0�011$1(1,1M1w1�1�1�1�1�1�1�1�1�122 2$2(2�2z3�3�3�56W6e6j6p6t6z6~6�6�6�6�6�6�6�6�6�6�6�6�6�6�6"7�7�7�7	88p8�8�8�8�8�8%9*949h9�9�9�9�9�9:
::Q:m:�:�:;y;�;�;�; <�<�<�<�<=4=;=C=H=L=P=y=�=�=�=�=�=�=�=�=�=�=*>0>4>8><>�>�>�>�>�>�>�>�>'?Y?`?d?h?l?p?t?x?|?�?�?�?�?�? � T   #0)0U0\0d0�0�0�0�011151�1�1B2�2�2'3A3J3R3q3{3�4�4�4�6�6�6�6~7�8�9�9x;�<   �   &0V0`0k0�2w3~3�3�3�3�3�3�3�3�3�3�3�3�3�3�34	4454J4p4�4�4�4�4�455@5�5�5�56'6s6�6�6�6�6�6�6�6�6�6�6�6�6�67777!7'7/767;7C7L7X7]7b7h7l7r7w7}7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�78$8<8X8�8�8�8�8�8�8H9N9T9Z9`9f9m9t9{9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9::::5:<:l:t:�:�:J=�=�=   |   F34�5�5�5�5�5"6*666�6�6�6�6�67�7�7�7 888�8�8�8�879?9G9S9_9�9�9�:�:!;);�;�;�<=�=�>�>�>�>??6???K?�?�?�?�?�?�?    �   000090�0�0�0�0�0�0�0�01 161A1[1f1n1~1�1�1�1�1�122&2Q2�2�2�2&3k3r3�3�3�34494]4�4�4�4�4�45+5P5[5j5�5�5�5�5666�7�7�7�788t8z8�8�8
99%9*9K9P9x9�9�9�9�9�9�9:�:�:;';~;=%=2=>=F=N=Z=�=�=�=�=�=>%>/>J>R>X>f>�>�>�>�>
?V?�?�?�?�?   �   060C0I011Z1l1{1q2w2�2�2�2�23M3�3�3�3�3�3�3�344'4R4m4t4}4�4�4�4�4�4�4�4�4555!5%5)5-5155595=5A5E5Z5�5D6�6�6�7�7�7�7�7�7�8�8�9�9�9�9 :::J:Q:[:m:�:�:�:�:�:�:�:�:�:;5;u;�;�;<<=Z=�=�=.>v>�>�?�? 0 �   30M0^0�0%1b1y1�2�243A3K3Y3b3l3�3�3�3�3�3�34F4{4�4�45d5�5�5g6s6�6�6�6�6�6�6�6777'7,7;7b7�7�7�7!8-8�8�8�8�8u9�9�:�:�;�=�? @ �   �011%1�1�1�1�1�12222-2\2b2j2�2�2�2�2�23333|3�3�34�4�4�4�455�5666$6)6:6B6H6R6X6b6h6r6{6�6�6�6�6�6�6�679!9'9f:m:R;�;<.<�<�<�<   P D   0�0A2�2�2�2�4�6�6�6�6�6�6�6�69�:�:�:�:�:=;F<�<�<L=�=�?�?�? ` `   	00$0T0�4�4�4�4�455/5A5S5e5w5�5�5�5�5�5�5�5E6�6�7(8K8�8S:�:�;�;�<d=�=>�>�>�>S?j?�?   p P   '01#1�1�2M3S3�3�34�4�4�4x558L8�;�;�;�;�;�;�;�;�;�;�;�;�;�<�<�<�<9=]=   � (   d7p9}9�9�9�9:�:
;�;�;�<�<?=�>�? � �   W0�0�0�0�0�1�1�1s2�2�233,3;3H3T3d3k3z3�3�3�3�3�3�3�34O4^4g4�4�4�4�46$6.9A9Y9y9�9�9:):V:�:�:�:�:�:�:;�;<E<f<o<�<�<�<�<�=�=�=�=1>�>�>�>�>�>Z?�?�?   � \   0N0X0(1e1o1�1�1�1
2�2�2�23"3B3b3�3�3�3�34"4B4b4�4�4�4�45"5B5b5�5�5�5�5�5�5�5�56 � �  1111 1$10141l1p1t1�1�1 22222222 2$2(2,2024282<2@2D2H2L2P2T2X2\2`2d2h2l2p2t2x2X3\3`3d3h3l3p3t3x3|3�3�3�3�3�3�3�3�3�3�3 44444444 4$4(4,404 555555�5�5�5�5�54686H6L6P6T6X6\6`6d6h6l6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�6�67 7$7(7,7074787<7@7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�8�8�8�8�8(9,9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9�9:p:t:x:|:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:�:;; � 4   ==$=,=4=<=D=L=T=\=d=l=t=|=�=�=�=�=�=�=�=�= � �   5555 5$5(5,5054585<5@5D5H5L5P5T5X5\5`5d5h5l5p5t5x5|5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5�5 66666666 6$6(6,6064686<6@6D6H6L6P6T6X6\6`6d6h6l6p6t6x6|6�6�6�6�6�6   � �  �4�4<5@5P5T5X5`5x5|5�5�5�5�5�5�5�5�5�5 666(6,60646<6T6d6h6x6|6�6�6�6�6�6�6�6�6�6�6�6�6�6�67$7(7,747L7\7`7t7x7|7�7�7�7�7�7�7�7�7�7�7�7 88 80848D8H8L8T8l8|8�8�8�8�8�8�8�8�8�8�8�8�8999(9,949L9\9`9p9t9x9�9�9�9�9�9�9�9�9�9�9�9�9:: :0:4:<:T:d:h:x:|:�:�:�:�:�:�:�:�:�:�:�: ;;;$;(;0;H;X;\;l;p;x;�;�;�;�;�;�;�;�;�;�; <<<$<4<8<H<L<P<X<p<�<�<�<�<�<�<�<�<�<�<�<�<�<�<�<= =$=4=8=H=L=T=l=|=�=�=�=�=�=�=L>T>\>`>h>|>�>�>�>�>�>�> ?$?0?8?X?|?�?�?�?�?�?�?     ,  0,080@0`0�0�0�0�0�0�0�0141@1H1h1�1�1�1�1�1�1�12<2H2P2p2�2�2�2�2�2�2 3 3D3P3X3x3�3�3�3�3�3 44(4L4X4`4�4�4�4�4�4�45505T5`5h5�5�5�5�5�566686\6h6p6�6�6�6�6�6�6�6�6�6�6�6�6�6�6 7707L7P7p7�7�7�7�7�7�7�788 8P8X8\8t8x8�8�8�8�8�8�8�8�8�8�89$9<9@9\9`9�9�9�9�9 : :<:@:\:`:�:�:�:�: ;;(;H;h;   �   0080P0h0�0�0�0�0�01,1L1t1�1�1�1�12,2H2`2|2�2�2�2�23<3�3�3�3�3�3�3�3�3�3�3�3�6�6�6�6�6�6�6�6�6�6 77777777 7$7(7,7074787<7@7D7H7L7P7T7X7\7`7d7h7l7p7t7x7|7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7�7 88888888 8$8(8,8084888�8�8�8�8�8�899999H=`>d>t>|>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>�>????$?,?4?<?D?L?T?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?�?   0     00@0H0                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                